configuration storage_routed_cfg of storage is
   for routed
   end for;
end storage_routed_cfg;
