library IEEE;
use IEEE.std_logic_1164.ALL;

entity counter4_tb is
end counter4_tb;

