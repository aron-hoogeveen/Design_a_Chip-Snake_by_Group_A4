configuration rng_synthesised_cfg of rng is
   for synthesised
   end for;
end rng_synthesised_cfg;
