library IEEE;
use IEEE.std_logic_1164.ALL;

entity shift_register_tb is
end shift_register_tb;

