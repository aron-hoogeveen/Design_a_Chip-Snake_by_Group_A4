library IEEE;
use IEEE.std_logic_1164.ALL;

entity snake_game_tb is
end snake_game_tb;

