library IEEE;
use IEEE.std_logic_1164.ALL;

entity storage_tb is
end storage_tb;

