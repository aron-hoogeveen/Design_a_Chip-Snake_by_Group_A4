configuration rng_tb_structural_cfg of rng_tb is
   for structural
      for all: rng use configuration work.rng_routed_cfg;
      end for;
   end for;
end rng_tb_structural_cfg;
