configuration storage_synthesised_cfg of storage is
   for synthesised
   end for;
end storage_synthesised_cfg;
