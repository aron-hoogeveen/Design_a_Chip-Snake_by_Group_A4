library IEEE;
use IEEE.std_logic_1164.ALL;

entity h_cnt_control_tb is
end h_cnt_control_tb;

