library IEEE;
use IEEE.std_logic_1164.ALL;

entity speed_tb is
end speed_tb;

