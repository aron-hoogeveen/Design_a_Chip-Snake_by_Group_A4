configuration mux_behaviour_cfg of mux is
   for behaviour
   end for;
end mux_behaviour_cfg;
