configuration rng_tb_behaviour_par of rng_tb is
   for behaviour
      for all: rng use configuration work.rng_routed_cfg;
      end for;
   end for;
end rng_tb_behaviour_par;
