library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

architecture structure of image_gen is
-- component decalaration
	component item_image is
   		port(clk   					: in  std_logic;
        		 reset 					: in  std_logic;
		  	  video_on   : in  std_logic;
       	 	 location_x : in  std_logic_vector(4 downto 0);
      	  	 location_y : in  std_logic_vector(4 downto 0);
     	   	 h_count    : in  std_logic_vector(8 downto 0);
    	    	 v_count    : in  std_logic_vector(9 downto 0);
   	     	 item      	: out std_logic);
	end component;

	component snake_image is
   		port(clk        : in  std_logic;
        		 reset      : in  std_logic;
        		 video_on   : in  std_logic;
        			loc_xL 				: in  std_logic_vector(4 downto 0);
		   	 loc_xH 				: in  std_logic_vector(4 downto 0);
        			loc_yL 				: in  std_logic_vector(4 downto 0);
		  	  loc_yH 				: in  std_logic_vector(4 downto 0);
        			h_count    : in  std_logic_vector(8 downto 0);
        			v_count    : in  std_logic_vector(9 downto 0);
        			snake      : out std_logic;
		  	  flag       : out std_logic);
	end component;

	component color_gen is
   	 port(clk      : in  std_logic;
     		  	reset    : in  std_logic;
     	    snake    : in  std_logic;
      	   item     : in  std_logic;
       	  video_on : in  std_logic;
        	 red      : out std_logic;
        	 green    : out std_logic;
        	 blue     : out std_logic);
	end component;

	signal snake_inter : std_logic;
	signal item_inter  : std_logic;

begin

item: item_image
	port map(clk   					=> clk,
        		  reset 					=> reset,
		  	   video_on   => video_on,
       	 	  location_x => item_x,
      	  	  location_y => item_y,
     	   	  h_count    => h_count,
    	    	  v_count    => v_count,
   	     	  item      	=> item_inter);

snake: snake_image
	port map(clk   			=> clk,
				reset 			=> reset,
        		 	video_on => video_on,
        				loc_xL 		=> snake_x_l,
		   	 	loc_xH 		=> snake_x_h,
        				loc_yL 		=> snake_y_l,
		  	  	loc_yH 		=> snake_y_h,
        				h_count  => h_count,
        				v_count  => v_count,
        				snake    => snake_inter,
		  	  	flag     => flag);

rgb: color_gen
	port map(clk      => clk,
      				reset    => reset,
        				snake    => snake_inter,
        				item     => item_inter,
        				video_on => video_on,
        				red      => red,
        				green    => green,
	         blue     => blue);

end structure;

