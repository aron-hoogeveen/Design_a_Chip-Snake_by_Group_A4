
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of storage is

  component CKND4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component LHD1BWP7T
    port(E, D : in std_logic; Q, QN : out std_logic);
  end component;

  component LND1BWP7T
    port(EN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(EN, D : in std_logic; Q : out std_logic);
  end component;

  component LHQD1BWP7T
    port(E, D : in std_logic; Q : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D4BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AN2D4BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component AN2D2BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component AOI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component TIELBWP7T
    port(ZN : out std_logic);
  end component;

  signal new_N : std_logic_vector(31 downto 0);
  signal new_corner_count : std_logic_vector(31 downto 0);
  signal new_state : std_logic_vector(4 downto 0);
  signal corner_count : std_logic_vector(31 downto 0);
  signal N : std_logic_vector(31 downto 0);
  signal state : std_logic_vector(4 downto 0);
  signal corner_check : std_logic_vector(5 downto 0);
  signal shift0 : std_logic_vector(5 downto 0);
  signal shift1 : std_logic_vector(5 downto 0);
  signal shift2 : std_logic_vector(5 downto 0);
  signal shift3 : std_logic_vector(5 downto 0);
  signal shift4 : std_logic_vector(5 downto 0);
  signal shift5 : std_logic_vector(5 downto 0);
  signal shift6 : std_logic_vector(5 downto 0);
  signal shift7 : std_logic_vector(5 downto 0);
  signal shift8 : std_logic_vector(5 downto 0);
  signal shift9 : std_logic_vector(5 downto 0);
  signal shift10 : std_logic_vector(5 downto 0);
  signal shift11 : std_logic_vector(5 downto 0);
  signal shift12 : std_logic_vector(5 downto 0);
  signal shift13 : std_logic_vector(5 downto 0);
  signal shift14 : std_logic_vector(5 downto 0);
  signal shift15 : std_logic_vector(5 downto 0);
  signal shift16 : std_logic_vector(5 downto 0);
  signal shift17 : std_logic_vector(5 downto 0);
  signal shift18 : std_logic_vector(5 downto 0);
  signal shift19 : std_logic_vector(5 downto 0);
  signal shift20 : std_logic_vector(5 downto 0);
  signal shift21 : std_logic_vector(5 downto 0);
  signal shift22 : std_logic_vector(5 downto 0);
  signal shift23 : std_logic_vector(5 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8 : std_logic;
  signal UNCONNECTED9, UNCONNECTED10, UNCONNECTED11, UNCONNECTED12, UNCONNECTED13 : std_logic;
  signal UNCONNECTED14, UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18 : std_logic;
  signal UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22, UNCONNECTED23 : std_logic;
  signal UNCONNECTED24, UNCONNECTED25, UNCONNECTED26, UNCONNECTED27, UNCONNECTED28 : std_logic;
  signal UNCONNECTED29, UNCONNECTED30, UNCONNECTED31, UNCONNECTED32, UNCONNECTED33 : std_logic;
  signal UNCONNECTED34, UNCONNECTED35, UNCONNECTED36, UNCONNECTED37, UNCONNECTED38 : std_logic;
  signal UNCONNECTED39, UNCONNECTED40, UNCONNECTED41, UNCONNECTED42, inc_add_286_38_n_0 : std_logic;
  signal inc_add_286_38_n_2, inc_add_286_38_n_4, inc_add_286_38_n_6, inc_add_286_38_n_8, inc_add_286_38_n_10 : std_logic;
  signal inc_add_286_38_n_12, inc_add_286_38_n_14, inc_add_286_38_n_16, inc_add_286_38_n_18, inc_add_286_38_n_20 : std_logic;
  signal inc_add_286_38_n_22, inc_add_286_38_n_24, inc_add_286_38_n_26, inc_add_286_38_n_28, inc_add_286_38_n_30 : std_logic;
  signal inc_add_286_38_n_32, inc_add_286_38_n_34, inc_add_286_38_n_36, inc_add_286_38_n_38, inc_add_286_38_n_40 : std_logic;
  signal inc_add_286_38_n_42, inc_add_286_38_n_44, inc_add_286_38_n_46, inc_add_286_38_n_48, inc_add_286_38_n_50 : std_logic;
  signal inc_add_286_38_n_52, inc_add_286_38_n_54, inc_add_286_38_n_56, inc_add_286_38_n_58, inc_add_1070_17_n_0 : std_logic;
  signal inc_add_1070_17_n_2, inc_add_1070_17_n_4, inc_add_1070_17_n_6, inc_add_1070_17_n_8, inc_add_1070_17_n_10 : std_logic;
  signal inc_add_1070_17_n_12, inc_add_1070_17_n_14, inc_add_1070_17_n_16, inc_add_1070_17_n_18, inc_add_1070_17_n_20 : std_logic;
  signal inc_add_1070_17_n_22, inc_add_1070_17_n_24, inc_add_1070_17_n_26, inc_add_1070_17_n_28, inc_add_1070_17_n_30 : std_logic;
  signal inc_add_1070_17_n_32, inc_add_1070_17_n_34, inc_add_1070_17_n_36, inc_add_1070_17_n_38, inc_add_1070_17_n_40 : std_logic;
  signal inc_add_1070_17_n_42, inc_add_1070_17_n_44, inc_add_1070_17_n_46, inc_add_1070_17_n_48, inc_add_1070_17_n_50 : std_logic;
  signal inc_add_1070_17_n_52, inc_add_1070_17_n_54, inc_add_1070_17_n_56, inc_add_1070_17_n_58, n_0 : std_logic;
  signal n_1, n_2, n_3, n_4, n_5 : std_logic;
  signal n_6, n_7, n_8, n_9, n_10 : std_logic;
  signal n_11, n_12, n_13, n_14, n_15 : std_logic;
  signal n_16, n_17, n_18, n_19, n_20 : std_logic;
  signal n_21, n_22, n_23, n_24, n_25 : std_logic;
  signal n_26, n_27, n_28, n_29, n_30 : std_logic;
  signal n_31, n_32, n_33, n_34, n_35 : std_logic;
  signal n_36, n_37, n_38, n_39, n_40 : std_logic;
  signal n_41, n_42, n_43, n_44, n_45 : std_logic;
  signal n_46, n_47, n_48, n_49, n_50 : std_logic;
  signal n_51, n_52, n_53, n_54, n_55 : std_logic;
  signal n_56, n_57, n_58, n_59, n_60 : std_logic;
  signal n_61, n_62, n_63, n_64, n_65 : std_logic;
  signal n_66, n_67, n_68, n_69, n_70 : std_logic;
  signal n_71, n_72, n_73, n_74, n_75 : std_logic;
  signal n_76, n_77, n_78, n_79, n_80 : std_logic;
  signal n_81, n_82, n_83, n_84, n_85 : std_logic;
  signal n_86, n_87, n_88, n_89, n_90 : std_logic;
  signal n_91, n_92, n_93, n_94, n_95 : std_logic;
  signal n_96, n_97, n_98, n_99, n_100 : std_logic;
  signal n_101, n_102, n_103, n_104, n_105 : std_logic;
  signal n_106, n_107, n_108, n_109, n_110 : std_logic;
  signal n_111, n_112, n_113, n_114, n_115 : std_logic;
  signal n_116, n_117, n_118, n_119, n_120 : std_logic;
  signal n_121, n_122, n_123, n_124, n_125 : std_logic;
  signal n_126, n_127, n_128, n_129, n_130 : std_logic;
  signal n_131, n_132, n_133, n_134, n_135 : std_logic;
  signal n_136, n_137, n_138, n_139, n_140 : std_logic;
  signal n_141, n_142, n_143, n_144, n_145 : std_logic;
  signal n_146, n_147, n_148, n_149, n_150 : std_logic;
  signal n_151, n_152, n_153, n_154, n_155 : std_logic;
  signal n_156, n_157, n_158, n_159, n_160 : std_logic;
  signal n_161, n_162, n_163, n_164, n_165 : std_logic;
  signal n_166, n_167, n_168, n_169, n_170 : std_logic;
  signal n_171, n_172, n_173, n_174, n_175 : std_logic;
  signal n_176, n_177, n_178, n_179, n_180 : std_logic;
  signal n_181, n_182, n_183, n_184, n_185 : std_logic;
  signal n_186, n_187, n_188, n_189, n_190 : std_logic;
  signal n_191, n_192, n_193, n_194, n_195 : std_logic;
  signal n_196, n_197, n_198, n_199, n_200 : std_logic;
  signal n_201, n_202, n_203, n_204, n_205 : std_logic;
  signal n_206, n_207, n_208, n_209, n_210 : std_logic;
  signal n_211, n_212, n_213, n_214, n_215 : std_logic;
  signal n_216, n_217, n_218, n_219, n_220 : std_logic;
  signal n_221, n_222, n_223, n_224, n_225 : std_logic;
  signal n_226, n_227, n_228, n_229, n_230 : std_logic;
  signal n_231, n_232, n_233, n_234, n_235 : std_logic;
  signal n_236, n_237, n_238, n_239, n_240 : std_logic;
  signal n_241, n_242, n_243, n_244, n_245 : std_logic;
  signal n_246, n_247, n_248, n_249, n_250 : std_logic;
  signal n_251, n_252, n_253, n_254, n_255 : std_logic;
  signal n_256, n_257, n_258, n_259, n_260 : std_logic;
  signal n_261, n_262, n_263, n_264, n_265 : std_logic;
  signal n_266, n_267, n_268, n_269, n_270 : std_logic;
  signal n_271, n_272, n_273, n_274, n_275 : std_logic;
  signal n_276, n_277, n_278, n_279, n_280 : std_logic;
  signal n_281, n_282, n_283, n_284, n_285 : std_logic;
  signal n_286, n_287, n_288, n_289, n_290 : std_logic;
  signal n_291, n_292, n_293, n_294, n_295 : std_logic;
  signal n_296, n_297, n_298, n_299, n_300 : std_logic;
  signal n_301, n_302, n_303, n_304, n_305 : std_logic;
  signal n_306, n_307, n_308, n_309, n_310 : std_logic;
  signal n_311, n_312, n_313, n_314, n_315 : std_logic;
  signal n_316, n_317, n_318, n_319, n_320 : std_logic;
  signal n_321, n_322, n_323, n_324, n_325 : std_logic;
  signal n_326, n_327, n_328, n_329, n_330 : std_logic;
  signal n_331, n_332, n_333, n_334, n_335 : std_logic;
  signal n_336, n_337, n_338, n_339, n_340 : std_logic;
  signal n_341, n_342, n_343, n_344, n_345 : std_logic;
  signal n_346, n_347, n_348, n_349, n_350 : std_logic;
  signal n_351, n_352, n_353, n_354, n_355 : std_logic;
  signal n_356, n_357, n_358, n_359, n_360 : std_logic;
  signal n_361, n_362, n_363, n_364, n_365 : std_logic;
  signal n_366, n_367, n_368, n_369, n_370 : std_logic;
  signal n_371, n_372, n_373, n_374, n_375 : std_logic;
  signal n_376, n_377, n_378, n_379, n_380 : std_logic;
  signal n_381, n_382, n_383, n_384, n_385 : std_logic;
  signal n_386, n_387, n_388, n_389, n_390 : std_logic;
  signal n_391, n_392, n_393, n_394, n_395 : std_logic;
  signal n_396, n_397, n_398, n_399, n_400 : std_logic;
  signal n_401, n_402, n_403, n_404, n_405 : std_logic;
  signal n_406, n_407, n_408, n_409, n_410 : std_logic;
  signal n_411, n_412, n_413, n_414, n_415 : std_logic;
  signal n_416, n_417, n_418, n_419, n_420 : std_logic;
  signal n_421, n_422, n_423, n_424, n_425 : std_logic;
  signal n_426, n_427, n_428, n_429, n_430 : std_logic;
  signal n_431, n_432, n_433, n_434, n_435 : std_logic;
  signal n_436, n_437, n_438, n_439, n_440 : std_logic;
  signal n_441, n_442, n_443, n_444, n_445 : std_logic;
  signal n_446, n_447, n_448, n_449, n_450 : std_logic;
  signal n_451, n_452, n_453, n_454, n_455 : std_logic;
  signal n_456, n_457, n_458, n_459, n_460 : std_logic;
  signal n_461, n_462, n_463, n_464, n_465 : std_logic;
  signal n_466, n_467, n_468, n_469, n_470 : std_logic;
  signal n_471, n_472, n_473, n_474, n_475 : std_logic;
  signal n_476, n_477, n_478, n_479, n_480 : std_logic;
  signal n_481, n_482, n_483, n_484, n_485 : std_logic;
  signal n_486, n_487, n_488, n_489, n_490 : std_logic;
  signal n_491, n_492, n_493, n_494, n_495 : std_logic;
  signal n_496, n_497, n_498, n_499, n_500 : std_logic;
  signal n_501, n_502, n_503, n_504, n_505 : std_logic;
  signal n_506, n_507, n_508, n_509, n_510 : std_logic;
  signal n_511, n_512, n_513, n_514, n_515 : std_logic;
  signal n_516, n_517, n_518, n_519, n_520 : std_logic;
  signal n_521, n_522, n_523, n_524, n_525 : std_logic;
  signal n_526, n_527, n_528, n_529, n_530 : std_logic;
  signal n_531, n_532, n_533, n_534, n_535 : std_logic;
  signal n_536, n_537, n_538, n_539, n_540 : std_logic;
  signal n_541, n_542, n_543, n_544, n_545 : std_logic;
  signal n_546, n_547, n_549, n_550, n_551 : std_logic;
  signal n_552, n_553, n_554, n_555, n_556 : std_logic;
  signal n_557, n_558, n_559, n_560, n_561 : std_logic;
  signal n_562, n_563, n_564, n_565, n_566 : std_logic;
  signal n_567, n_568, n_569, n_570, n_571 : std_logic;
  signal n_572, n_573, n_574, n_575, n_576 : std_logic;
  signal n_577, n_578, n_579, n_580, n_581 : std_logic;
  signal n_582, n_583, n_584, n_585, n_586 : std_logic;
  signal n_587, n_588, n_589, n_590, n_591 : std_logic;
  signal n_592, n_593, n_594, n_595, n_596 : std_logic;
  signal n_597, n_598, n_599, n_600, n_601 : std_logic;
  signal n_602, n_603, n_604, n_605, n_606 : std_logic;
  signal n_607, n_608, n_609, n_610, n_611 : std_logic;
  signal n_612, n_613, n_614, n_615, n_616 : std_logic;
  signal n_617, n_618, n_619, n_620, n_621 : std_logic;
  signal n_622, n_623, n_624, n_625, n_626 : std_logic;
  signal n_627, n_628, n_629, n_630, n_631 : std_logic;
  signal n_632, n_633, n_634, n_635, n_636 : std_logic;
  signal n_637, n_638, n_639, n_640, n_641 : std_logic;
  signal n_642, n_643, n_644, n_645, n_646 : std_logic;
  signal n_647, n_648, n_649, n_650, n_651 : std_logic;
  signal n_652, n_653, n_654, n_655, n_656 : std_logic;
  signal n_657, n_658, n_659, n_660, n_661 : std_logic;
  signal n_662, n_663, n_664, n_665, n_666 : std_logic;
  signal n_667, n_668, n_669, n_670, n_671 : std_logic;
  signal n_672, n_673, n_674, n_675, n_676 : std_logic;
  signal n_677, n_678, n_679, n_680, n_681 : std_logic;
  signal n_682, n_683, n_684, n_685, n_686 : std_logic;
  signal n_687, n_688, n_689, n_690, n_691 : std_logic;
  signal n_692, n_693, n_694, n_695, n_696 : std_logic;
  signal n_697, n_698, n_699, n_700, n_701 : std_logic;
  signal n_702, n_703, n_704, n_705, n_706 : std_logic;
  signal n_707, n_708, n_709, n_710, n_711 : std_logic;
  signal n_712, n_713, n_714, n_715, n_716 : std_logic;
  signal n_717, n_718, n_719, n_720, n_721 : std_logic;
  signal n_722, n_723, n_724, n_725, n_726 : std_logic;
  signal n_727, n_728, n_729, n_730, n_731 : std_logic;
  signal n_732, n_733, n_734, n_735, n_736 : std_logic;
  signal n_737, n_738, n_739, n_740, n_741 : std_logic;
  signal n_742, n_743, n_744, n_745, n_746 : std_logic;
  signal n_747, n_748, n_749, n_750, n_751 : std_logic;
  signal n_752, n_753, n_754, n_755, n_756 : std_logic;
  signal n_757, n_758, n_759, n_760, n_761 : std_logic;
  signal n_762, n_763, n_764, n_765, n_766 : std_logic;
  signal n_767, n_768, n_769, n_770, n_771 : std_logic;
  signal n_772, n_773, n_774, n_775, n_776 : std_logic;
  signal n_777, n_778, n_779, n_780, n_781 : std_logic;
  signal n_782, n_783, n_784, n_785, n_786 : std_logic;
  signal n_787, n_788, n_789, n_790, n_791 : std_logic;
  signal n_792, n_793, n_794, n_795, n_796 : std_logic;
  signal n_797, n_798, n_799, n_800, n_801 : std_logic;
  signal n_802, n_803, n_804, n_805, n_806 : std_logic;
  signal n_807, n_808, n_809, n_810, n_811 : std_logic;
  signal n_812, n_813, n_814, n_815, n_816 : std_logic;
  signal n_817, n_818, n_819, n_820, n_821 : std_logic;
  signal n_822, n_823, n_824, n_825, n_826 : std_logic;
  signal n_827, n_828, n_829, n_830, n_831 : std_logic;
  signal n_832, n_833, n_834, n_835, n_836 : std_logic;
  signal n_837, n_838, n_839, n_840, n_841 : std_logic;
  signal n_842, n_843, n_844, n_845, n_846 : std_logic;
  signal n_847, n_848, n_849, n_850, n_851 : std_logic;
  signal n_852, n_853, n_854, n_855, n_856 : std_logic;
  signal n_857, n_858, n_859, n_860, n_861 : std_logic;
  signal n_862, n_863, n_864, n_865, n_866 : std_logic;
  signal n_867, n_868, n_869, n_870, n_871 : std_logic;
  signal n_872, n_873, n_874, n_875, n_876 : std_logic;
  signal n_877, n_878, n_879, n_880, n_881 : std_logic;
  signal n_882, n_883, n_884, n_885, n_886 : std_logic;
  signal n_887, n_888, n_889, n_890, n_891 : std_logic;
  signal n_892, n_893, n_894, n_895, n_896 : std_logic;
  signal n_897, n_898, n_899, n_900, n_901 : std_logic;
  signal n_902, n_903, n_904, n_905, n_906 : std_logic;
  signal n_907, n_908, n_909, n_910, n_911 : std_logic;
  signal n_912, n_913, n_914, n_915, n_916 : std_logic;
  signal n_917, n_918, n_919, n_920, n_921 : std_logic;
  signal n_922, n_923, n_924, n_925, n_926 : std_logic;
  signal n_927, n_928, n_929, n_930, n_931 : std_logic;
  signal n_932, n_933, n_934, n_935, n_936 : std_logic;
  signal n_937, n_938, n_939, n_940, n_941 : std_logic;
  signal n_942, n_943, n_944, n_945, n_946 : std_logic;
  signal n_947, n_948, n_949, n_950, n_951 : std_logic;
  signal n_952, n_953, n_954, n_955, n_956 : std_logic;
  signal n_957, n_958, n_959, n_960, n_961 : std_logic;
  signal n_962, n_963, n_964, n_965, n_966 : std_logic;
  signal n_967, n_968, n_969, n_970, n_971 : std_logic;
  signal n_972, n_973, n_974, n_975, n_976 : std_logic;
  signal n_977, n_978, n_979, n_980, n_981 : std_logic;
  signal n_982, n_983, n_984, n_985, n_986 : std_logic;
  signal n_987, n_988, n_989, n_990, n_991 : std_logic;
  signal n_992, n_993, n_994, n_995, n_996 : std_logic;
  signal n_997, n_998, n_999, n_1000, n_1001 : std_logic;
  signal n_1002, n_1003, n_1004, n_1005, n_1006 : std_logic;
  signal n_1007, n_1008, n_1009, n_1010, n_1011 : std_logic;
  signal n_1012, n_1013, n_1014, n_1015, n_1016 : std_logic;
  signal n_1017, n_1018, n_1019, n_1020, n_1021 : std_logic;
  signal n_1022, n_1023, n_1024, n_1025, n_1026 : std_logic;
  signal n_1027, n_1028, n_1029, n_1030, n_1031 : std_logic;
  signal n_1032, n_1033, n_1034, n_1035, n_1036 : std_logic;
  signal n_1037, n_1038, n_1039, n_1040, n_1041 : std_logic;
  signal n_1042, n_1043, n_1044, n_1045, n_1046 : std_logic;
  signal n_1047, n_1048, n_1049, n_1050, n_1051 : std_logic;
  signal n_1052, n_1053, n_1054, n_1055, n_1056 : std_logic;
  signal n_1057, n_1058, n_1059, n_1060, n_1061 : std_logic;
  signal n_1062, n_1063, n_1064, n_1065, n_1066 : std_logic;
  signal n_1067, n_1068, n_1069, n_1070, n_1071 : std_logic;
  signal n_1072, n_1073, n_1074, n_1075, n_1076 : std_logic;
  signal n_1077, n_1078, n_1079, n_1080, n_1081 : std_logic;
  signal n_1082, n_1083, n_1084, n_1085, n_1086 : std_logic;
  signal n_1087, n_1088, n_1089, n_1090, n_1091 : std_logic;
  signal n_1092, n_1093, n_1094, n_1095, n_1096 : std_logic;
  signal n_1097, n_1098, n_1099, n_1100, n_1101 : std_logic;
  signal n_1102, n_1103, n_1104, n_1105, n_1106 : std_logic;
  signal n_1107, n_1108, n_1109, n_1110, n_1111 : std_logic;
  signal n_1112, n_1113, n_1114, n_1115, n_1116 : std_logic;
  signal n_1117, n_1118, n_1119, n_1120, n_1121 : std_logic;
  signal n_1122, n_1123, n_1124, n_1125, n_1126 : std_logic;
  signal n_1127, n_1128, n_1129, n_1130, n_1131 : std_logic;
  signal n_1132, n_1133, n_1134, n_1135, n_1136 : std_logic;
  signal n_1137, n_1138, n_1139, n_1140, n_1141 : std_logic;
  signal n_1142, n_1143, n_1144, n_1145, n_1146 : std_logic;
  signal n_1147, n_1148, n_1149, n_1150, n_1151 : std_logic;
  signal n_1152, n_1153, n_1154, n_1155, n_1156 : std_logic;
  signal n_1157, n_1158, n_1159, n_1160, n_1161 : std_logic;
  signal n_1162, n_1163, n_1164, n_1165, n_1166 : std_logic;
  signal n_1167, n_1168, n_1169, n_1170, n_1171 : std_logic;
  signal n_1172, n_1173, n_1174, n_1175, n_1176 : std_logic;
  signal n_1177, n_1178, n_1179, n_1180, n_1181 : std_logic;
  signal n_1182, n_1183, n_1184, n_1185, n_1186 : std_logic;
  signal n_1187, n_1188, n_1189, n_1190, n_1191 : std_logic;
  signal n_1192, n_1193, n_1194, n_1195, n_1196 : std_logic;
  signal n_1197, n_1198, n_1199, n_1200, n_1201 : std_logic;
  signal n_1202, n_1203, n_1204, n_1205, n_1206 : std_logic;
  signal n_1207, n_1208, n_1209, n_1210, n_1211 : std_logic;
  signal n_1212, n_1214, n_1215, n_1216, n_1217 : std_logic;
  signal n_1218, n_1219, n_1220, n_1221, n_1222 : std_logic;
  signal n_1223, n_1224, n_1225, n_1226, n_1227 : std_logic;
  signal n_1228, n_1229, n_1230, n_1231, n_1232 : std_logic;
  signal n_1233, n_1234, n_1235, n_1236, n_1237 : std_logic;
  signal n_1238, n_1239, n_1240, n_1241, n_1242 : std_logic;
  signal n_1243, n_1244, n_1245, n_1246, n_1247 : std_logic;
  signal n_1248, n_1249, n_1250, n_1251, n_1252 : std_logic;
  signal n_1253, n_1254, n_1255, n_1256, n_1257 : std_logic;
  signal n_1258, n_1259, n_1260, n_1261, n_1262 : std_logic;
  signal n_1263, n_1264, n_1265, n_1266, n_1267 : std_logic;
  signal n_1268, n_1269, n_1270, n_1271, n_1272 : std_logic;
  signal n_1273, n_1274, n_1275, n_1276, n_1277 : std_logic;
  signal n_1278, n_1279, n_1280, n_1281, n_1282 : std_logic;
  signal n_1283, n_1284, n_1285, n_1286, n_1287 : std_logic;
  signal n_1288, n_1289, n_1290, n_1291, n_1292 : std_logic;
  signal n_1293, n_1294, n_1295, n_1296, n_1297 : std_logic;
  signal n_1298, n_1299, n_1300, n_1301, n_1302 : std_logic;
  signal n_1303, n_1304, n_1305, n_1306, n_1307 : std_logic;
  signal n_1309, n_1310, n_1311, n_1312, n_1313 : std_logic;
  signal n_1314, n_1315, n_1316, n_1317, n_1318 : std_logic;
  signal n_1319, n_1320, n_1321, n_1322, n_1323 : std_logic;
  signal n_1324, n_1325, n_1326, n_1327, n_1328 : std_logic;
  signal n_1329, n_1330, n_1331, n_1332, n_1333 : std_logic;
  signal n_1334, n_1335, n_1336, n_1337, n_1338 : std_logic;
  signal n_1339, n_1340, n_1341, n_1342, n_1343 : std_logic;
  signal n_1344, n_1345, n_1346, n_1347, n_1348 : std_logic;
  signal n_1349, n_1350, n_1351, n_1352, n_1353 : std_logic;
  signal n_1354, n_1355, n_1357, n_1358, n_1359 : std_logic;
  signal n_1360, n_1361, n_1362, n_1363, n_1364 : std_logic;
  signal n_1365, n_1366, n_1367, n_1368, n_1369 : std_logic;
  signal n_1370, n_1371, n_1372, n_1373, n_1374 : std_logic;
  signal n_1375, n_1376, n_1377, n_1378, n_1379 : std_logic;
  signal n_1380, n_1381, n_1382, n_1383, n_1384 : std_logic;
  signal n_1385, n_1386, n_1387, n_1388, n_1389 : std_logic;
  signal n_1390, n_1391, n_1392, n_1393, n_1394 : std_logic;
  signal n_1395, n_1396, n_1397, n_1399, n_1400 : std_logic;
  signal n_1401, n_1402, n_1403, n_1404, n_1405 : std_logic;
  signal n_1406, n_1407, n_1408, n_1409, n_1410 : std_logic;
  signal n_1411, n_1413, n_1414, n_1415, n_1416 : std_logic;
  signal n_1417, n_1418, n_1419, n_1420, n_1421 : std_logic;
  signal n_1422, n_1423, n_1424, n_1425, n_1426 : std_logic;
  signal n_1564, n_1565, n_1566, n_1567, n_1568 : std_logic;
  signal n_1569, n_1570, n_1571, n_1572, n_1573 : std_logic;
  signal n_1574, n_1575, n_1578, n_1579, n_1580 : std_logic;
  signal n_1581, n_1582, n_1583, n_1584, n_1585 : std_logic;
  signal n_1587, n_1588, n_1589, n_1590, n_1591 : std_logic;
  signal n_1592, n_1593, n_1594, n_1595, n_1596 : std_logic;
  signal n_1597, n_1598, n_1599, n_1600, n_1601 : std_logic;
  signal n_1602, n_1603, n_1604, n_1605, n_1606 : std_logic;
  signal n_1607, n_1608, n_1609, n_1610, n_1611 : std_logic;
  signal n_1612, n_1613, n_1614, n_1615, n_1616 : std_logic;
  signal n_1617, n_1618, n_1619, n_1620, n_1621 : std_logic;
  signal n_1622, n_1623, n_1624, n_1625, n_1626 : std_logic;
  signal n_1627, n_1628, n_1629, n_1630, n_1631 : std_logic;
  signal n_1632, n_1633, n_1634, n_1635, n_1636 : std_logic;
  signal n_1637, n_1638, n_1639, n_1640, n_1641 : std_logic;
  signal n_1642, n_1643, n_1644, n_1645, n_1646 : std_logic;
  signal n_1647, n_1648, n_1649, n_1650, n_1651 : std_logic;
  signal n_1652, n_1653, n_1654, n_1657, n_1662 : std_logic;
  signal n_1663, n_1670, n_1671, n_1672, n_1673 : std_logic;
  signal n_1674, n_1675, n_1676, n_1677, n_1678 : std_logic;
  signal n_1679, n_1680, n_1681, n_1682, n_1683 : std_logic;
  signal n_1684, n_1685, n_1686, n_1687, n_1688 : std_logic;
  signal n_1689, n_1690, n_1691, n_1692, n_1693 : std_logic;
  signal n_1694, n_1695, n_1696, n_1697, n_1698 : std_logic;
  signal n_1699, n_1700, n_1701, n_1703, n_1704 : std_logic;
  signal n_1705, n_1718, n_1731, n_1732, n_1733 : std_logic;
  signal n_1734, n_1735, n_1736, n_1737, n_1738 : std_logic;
  signal n_1739, n_1740, n_1742, n_1747, n_1748 : std_logic;
  signal n_1749, sub_868_22_n_0, sub_868_22_n_2, sub_868_22_n_4, sub_868_22_n_6 : std_logic;
  signal sub_868_22_n_8, sub_868_22_n_10, sub_868_22_n_12, sub_868_22_n_14, sub_868_22_n_16 : std_logic;
  signal sub_868_22_n_18, sub_868_22_n_20, sub_868_22_n_22, sub_868_22_n_24, sub_868_22_n_26 : std_logic;
  signal sub_868_22_n_28, sub_868_22_n_30, sub_868_22_n_32, sub_868_22_n_34, sub_868_22_n_36 : std_logic;
  signal sub_868_22_n_38, sub_868_22_n_40, sub_868_22_n_42, sub_868_22_n_44, sub_868_22_n_46 : std_logic;
  signal sub_868_22_n_48, sub_868_22_n_50, sub_868_22_n_52, sub_868_22_n_54, sub_868_22_n_56 : std_logic;
  signal sub_868_22_n_58 : std_logic;

begin

  send_new_corner_clear <= audio(7);
  item_send_flag <= audio(7);
  head_send_flag <= audio(7);
  remove_item_clear <= audio(7);
  audio(0) <= audio(7);
  audio(1) <= audio(7);
  audio(2) <= audio(7);
  audio(3) <= audio(7);
  audio(4) <= audio(7);
  audio(5) <= audio(7);
  audio(6) <= audio(7);
  g7522 : CKND4BWP7T port map(I => n_1651, ZN => snake_send_flag);
  H_S_reg_0_0 : LHD1BWP7T port map(E => n_1353, D => n_1312, Q => UNCONNECTED, QN => n_1350);
  H_S_reg_0_1 : LHD1BWP7T port map(E => n_1353, D => n_1311, Q => UNCONNECTED0, QN => n_1346);
  H_S_reg_0_2 : LHD1BWP7T port map(E => n_1353, D => n_1310, Q => UNCONNECTED1, QN => n_1347);
  H_S_reg_0_3 : LHD1BWP7T port map(E => n_1353, D => n_1309, Q => UNCONNECTED2, QN => n_1354);
  H_S_reg_0_4 : LHD1BWP7T port map(E => n_1353, D => n_1313, Q => UNCONNECTED3, QN => n_1351);
  H_S_reg_0_5 : LHD1BWP7T port map(E => n_1353, D => n_1315, Q => UNCONNECTED4, QN => n_1352);
  H_S_reg_0_6 : LHD1BWP7T port map(E => n_1353, D => n_1314, Q => UNCONNECTED5, QN => n_1337);
  H_S_reg_0_7 : LHD1BWP7T port map(E => n_1353, D => n_1291, Q => UNCONNECTED6, QN => n_1343);
  H_S_reg_0_8 : LHD1BWP7T port map(E => n_1353, D => n_1292, Q => UNCONNECTED7, QN => n_1348);
  H_S_reg_0_9 : LHD1BWP7T port map(E => n_1353, D => n_1317, Q => UNCONNECTED8, QN => n_1344);
  H_S_reg_0_10 : LHD1BWP7T port map(E => n_1353, D => n_1300, Q => UNCONNECTED9, QN => n_1345);
  H_S_reg_0_11 : LHD1BWP7T port map(E => n_1353, D => n_1293, Q => UNCONNECTED10, QN => n_1349);
  I_S_reg_0_0 : LHD1BWP7T port map(E => n_1386, D => n_1301, Q => UNCONNECTED11, QN => n_1366);
  I_S_reg_0_1 : LHD1BWP7T port map(E => n_1386, D => n_1299, Q => UNCONNECTED12, QN => n_1370);
  I_S_reg_0_2 : LHD1BWP7T port map(E => n_1386, D => n_1319, Q => UNCONNECTED13, QN => n_1374);
  I_S_reg_0_3 : LHD1BWP7T port map(E => n_1386, D => n_1298, Q => UNCONNECTED14, QN => n_1376);
  I_S_reg_0_4 : LHD1BWP7T port map(E => n_1386, D => n_1297, Q => UNCONNECTED15, QN => n_1380);
  I_S_reg_0_5 : LHD1BWP7T port map(E => n_1386, D => n_1296, Q => UNCONNECTED16, QN => n_1388);
  I_S_reg_0_6 : LHD1BWP7T port map(E => n_1386, D => n_1316, Q => UNCONNECTED17, QN => n_1365);
  I_S_reg_0_7 : LHD1BWP7T port map(E => n_1386, D => n_1295, Q => UNCONNECTED18, QN => n_1371);
  I_S_reg_0_8 : LHD1BWP7T port map(E => n_1386, D => n_1294, Q => UNCONNECTED19, QN => n_1377);
  I_S_reg_0_9 : LHD1BWP7T port map(E => n_1386, D => n_1302, Q => UNCONNECTED20, QN => n_1382);
  I_S_reg_0_10 : LHD1BWP7T port map(E => n_1386, D => n_1327, Q => UNCONNECTED21, QN => n_1368);
  I_S_reg_0_11 : LHD1BWP7T port map(E => n_1386, D => n_1330, Q => UNCONNECTED22, QN => n_1385);
  I_S_reg_1_0 : LND1BWP7T port map(EN => n_1384, D => n_1331, Q => UNCONNECTED23, QN => n_1367);
  I_S_reg_1_1 : LND1BWP7T port map(EN => n_1384, D => n_1329, Q => UNCONNECTED24, QN => n_1369);
  I_S_reg_1_2 : LND1BWP7T port map(EN => n_1384, D => n_1328, Q => UNCONNECTED25, QN => n_1372);
  I_S_reg_1_3 : LND1BWP7T port map(EN => n_1384, D => n_1318, Q => UNCONNECTED26, QN => n_1373);
  I_S_reg_1_4 : LND1BWP7T port map(EN => n_1384, D => n_1326, Q => UNCONNECTED27, QN => n_1375);
  I_S_reg_1_5 : LND1BWP7T port map(EN => n_1384, D => n_1325, Q => UNCONNECTED28, QN => n_1378);
  I_S_reg_1_6 : LND1BWP7T port map(EN => n_1384, D => n_1324, Q => UNCONNECTED29, QN => n_1379);
  I_S_reg_1_7 : LND1BWP7T port map(EN => n_1384, D => n_1332, Q => UNCONNECTED30, QN => n_1381);
  I_S_reg_1_8 : LND1BWP7T port map(EN => n_1384, D => n_1323, Q => UNCONNECTED31, QN => n_1383);
  I_S_reg_1_9 : LND1BWP7T port map(EN => n_1384, D => n_1322, Q => UNCONNECTED32, QN => n_1387);
  I_S_reg_1_10 : LND1BWP7T port map(EN => n_1384, D => n_1321, Q => UNCONNECTED33, QN => n_1363);
  I_S_reg_1_11 : LND1BWP7T port map(EN => n_1384, D => n_1320, Q => UNCONNECTED34, QN => n_1364);
  S_S_reg_0_0 : LND1BWP7T port map(EN => n_1401, D => n_1341, Q => UNCONNECTED35, QN => n_1400);
  S_S_reg_0_1 : LND1BWP7T port map(EN => n_1401, D => n_1360, Q => UNCONNECTED36, QN => n_1395);
  S_S_reg_0_2 : LND1BWP7T port map(EN => n_1401, D => n_1359, Q => UNCONNECTED37, QN => n_155);
  S_S_reg_0_3 : LND1BWP7T port map(EN => n_1401, D => n_1358, Q => UNCONNECTED38, QN => n_1402);
  S_S_reg_0_4 : LND1BWP7T port map(EN => n_1401, D => n_1357, Q => UNCONNECTED39, QN => n_1394);
  S_S_reg_0_5 : LND1BWP7T port map(EN => n_1401, D => n_1335, Q => UNCONNECTED40, QN => n_1399);
  new_N_reg_0 : LNQD1BWP7T port map(EN => n_1651, D => n_152, Q => new_N(0));
  new_corner_count_reg_0 : LHQD1BWP7T port map(E => n_1657, D => n_146, Q => new_corner_count(0));
  new_state_reg_2 : LHQD1BWP7T port map(E => n_1649, D => n_1415, Q => new_state(2));
  new_state_reg_3 : LHQD1BWP7T port map(E => n_1649, D => n_1414, Q => new_state(3));
  new_state_reg_4 : LHQD1BWP7T port map(E => n_1649, D => n_1420, Q => new_state(4));
  snake_list_reg_0 : LHD1BWP7T port map(E => n_1652, D => n_1411, Q => UNCONNECTED41, QN => n_1417);
  tail_reg : LHD1BWP7T port map(E => n_1651, D => n_1404, Q => UNCONNECTED42, QN => n_1407);
  g12536 : IND4D0BWP7T port map(A1 => n_1569, B1 => n_1279, B2 => n_1307, B3 => n_1426, ZN => n_1649);
  g12537 : NR4D0BWP7T port map(A1 => n_1425, A2 => n_1410, A3 => n_1579, A4 => n_1734, ZN => n_1426);
  g12538 : AO21D0BWP7T port map(A1 => n_1274, A2 => n_1209, B => n_1571, Z => n_1425);
  g12539 : AN2D1BWP7T port map(A1 => n_1650, A2 => n_1654, Z => n_1571);
  g12540 : IND4D0BWP7T port map(A1 => corner_count(8), B1 => n_1212, B2 => corner_count(0), B3 => n_1424, ZN => n_1650);
  g12541 : INR4D0BWP7T port map(A1 => n_1423, B1 => corner_count(9), B2 => corner_count(12), B3 => corner_count(10), ZN => n_1424);
  g12542 : INR4D0BWP7T port map(A1 => n_1422, B1 => corner_count(13), B2 => corner_count(16), B3 => corner_count(14), ZN => n_1423);
  g12543 : INR4D0BWP7T port map(A1 => n_1421, B1 => corner_count(17), B2 => corner_count(20), B3 => corner_count(18), ZN => n_1422);
  g12544 : INR4D0BWP7T port map(A1 => n_1419, B1 => corner_count(21), B2 => corner_count(5), B3 => corner_count(4), ZN => n_1421);
  g12545 : AN4D1BWP7T port map(A1 => n_1418, A2 => n_1277, A3 => n_1279, A4 => n_1203, Z => n_1420);
  g12546 : INR4D0BWP7T port map(A1 => n_1416, B1 => corner_count(6), B2 => corner_count(7), B3 => corner_count(3), ZN => n_1419);
  g12547 : NR4D0BWP7T port map(A1 => n_1749, A2 => n_1303, A3 => new_item_clear, A4 => clear_corner_flag, ZN => n_1418);
  g12549 : INVD4BWP7T port map(I => n_1417, ZN => snake_list(0));
  g12550 : INR4D0BWP7T port map(A1 => n_1408, B1 => corner_count(11), B2 => corner_count(19), B3 => corner_count(15), ZN => n_1416);
  g12551 : IND3D0BWP7T port map(A1 => n_1733, B1 => n_1409, B2 => n_1342, ZN => n_1415);
  g12552 : OR4D0BWP7T port map(A1 => n_1406, A2 => n_1734, A3 => n_1303, A4 => n_1568, Z => n_1414);
  g12553 : ND2D0BWP7T port map(A1 => n_1413, A2 => n_1279, ZN => n_1652);
  g12554 : NR2D0BWP7T port map(A1 => n_1410, A2 => n_1654, ZN => n_1413);
  g12556 : INR2D0BWP7T port map(A1 => tail, B1 => n_1651, ZN => n_1411);
  g12557 : AOI211D0BWP7T port map(A1 => n_1572, A2 => n_1747, B => n_1334, C => n_1403, ZN => n_1409);
  g12558 : IND4D0BWP7T port map(A1 => n_1572, B1 => n_1222, B2 => n_1276, B3 => n_1396, ZN => n_1410);
  g12559 : INR4D0BWP7T port map(A1 => n_1393, B1 => corner_count(22), B2 => corner_count(24), B3 => corner_count(23), ZN => n_1408);
  g12561 : INVD4BWP7T port map(I => n_1407, ZN => tail);
  g12562 : IND2D0BWP7T port map(A1 => n_1567, B1 => n_1392, ZN => n_1406);
  g12563 : OA221D0BWP7T port map(A1 => n_1283, A2 => n_1573, B1 => n_1397, B2 => n_1651, C => n_1336, Z => n_1405);
  g12564 : AN2D1BWP7T port map(A1 => n_1737, A2 => n_1397, Z => n_1566);
  g12565 : AN2D1BWP7T port map(A1 => n_1653, A2 => n_1397, Z => n_1567);
  g12566 : IAO21D0BWP7T port map(A1 => n_1569, A2 => n_1733, B => n_1397, ZN => n_1404);
  g12567 : OA21D0BWP7T port map(A1 => n_1737, A2 => n_1732, B => n_1397, Z => n_1403);
  g12569 : INVD4BWP7T port map(I => n_1402, ZN => snake_output0(3));
  g12571 : INVD4BWP7T port map(I => n_1400, ZN => snake_output0(0));
  g12573 : INVD4BWP7T port map(I => n_1399, ZN => snake_output0(5));
  g12575 : INVD4BWP7T port map(I => n_155, ZN => snake_output0(2));
  g12576 : NR4D0BWP7T port map(A1 => n_1391, A2 => n_1568, A3 => n_1303, A4 => n_1305, ZN => n_1396);
  g12578 : INVD4BWP7T port map(I => n_1395, ZN => snake_output0(1));
  g12580 : INVD4BWP7T port map(I => n_1394, ZN => snake_output0(4));
  g12581 : ND4D0BWP7T port map(A1 => n_1389, A2 => n_1390, A3 => n_1262, A4 => n_1215, ZN => n_1397);
  g12582 : NR4D0BWP7T port map(A1 => n_1361, A2 => corner_count(26), A3 => corner_count(25), A4 => corner_count(27), ZN => n_1393);
  g12583 : AOI32D0BWP7T port map(A1 => n_1572, A2 => n_1585, A3 => n_1273, B1 => n_1306, B2 => send_corner_flag, ZN => n_1392);
  g12584 : AOI211D0BWP7T port map(A1 => n_1362, A2 => n_1305, B => n_1278, C => n_1739, ZN => n_1401);
  g12585 : IIND4D0BWP7T port map(A1 => n_1663, A2 => new_item_clear, B1 => n_1287, B2 => n_1275, ZN => n_1391);
  g12586 : NR4D0BWP7T port map(A1 => n_1355, A2 => n_1284, A3 => n_1246, A4 => n_1244, ZN => n_1390);
  g12587 : NR4D0BWP7T port map(A1 => n_1338, A2 => n_1285, A3 => n_1289, A4 => n_1249, ZN => n_1389);
  g12589 : INVD4BWP7T port map(I => n_1388, ZN => item_out_food(5));
  g12591 : INVD4BWP7T port map(I => n_1387, ZN => item_out_power_up(9));
  g12593 : INVD4BWP7T port map(I => n_1385, ZN => item_out_food(11));
  g12595 : INVD4BWP7T port map(I => n_1383, ZN => item_out_power_up(8));
  g12597 : INVD4BWP7T port map(I => n_1382, ZN => item_out_food(9));
  g12599 : INVD4BWP7T port map(I => n_1381, ZN => item_out_power_up(7));
  g12601 : INVD4BWP7T port map(I => n_1380, ZN => item_out_food(4));
  g12603 : INVD4BWP7T port map(I => n_1379, ZN => item_out_power_up(6));
  g12605 : INVD4BWP7T port map(I => n_1378, ZN => item_out_power_up(5));
  g12607 : INVD4BWP7T port map(I => n_1377, ZN => item_out_food(8));
  g12609 : INVD4BWP7T port map(I => n_1376, ZN => item_out_food(3));
  g12611 : INVD4BWP7T port map(I => n_1375, ZN => item_out_power_up(4));
  g12613 : INVD4BWP7T port map(I => n_1374, ZN => item_out_food(2));
  g12615 : INVD4BWP7T port map(I => n_1373, ZN => item_out_power_up(3));
  g12617 : INVD4BWP7T port map(I => n_1372, ZN => item_out_power_up(2));
  g12619 : INVD4BWP7T port map(I => n_1371, ZN => item_out_food(7));
  g12621 : INVD4BWP7T port map(I => n_1370, ZN => item_out_food(1));
  g12623 : INVD4BWP7T port map(I => n_1369, ZN => item_out_power_up(1));
  g12625 : INVD4BWP7T port map(I => n_1368, ZN => item_out_food(10));
  g12627 : INVD4BWP7T port map(I => n_1367, ZN => item_out_power_up(0));
  g12629 : INVD4BWP7T port map(I => n_1366, ZN => item_out_food(0));
  g12631 : INVD4BWP7T port map(I => n_1365, ZN => item_out_food(6));
  g12633 : INVD4BWP7T port map(I => n_1364, ZN => item_out_power_up(11));
  g12635 : INVD4BWP7T port map(I => n_1363, ZN => item_out_power_up(10));
  g12636 : INR2D0BWP7T port map(A1 => n_1580, B1 => n_1339, ZN => n_1362);
  g12637 : IND2D0BWP7T port map(A1 => corner_count(28), B1 => n_1340, ZN => n_1361);
  g12638 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(1), B1 => n_1670, B2 => new_tail(1), C => n_1739, Z => n_1360);
  g12639 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(2), B1 => n_1670, B2 => new_tail(2), C => n_1739, Z => n_1359);
  g12640 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(3), B1 => n_1670, B2 => new_tail(3), C => n_1739, Z => n_1358);
  g12641 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(4), B1 => n_1670, B2 => new_tail(4), C => n_1739, Z => n_1357);
  g12643 : ND4D0BWP7T port map(A1 => n_1288, A2 => n_1290, A3 => n_1234, A4 => n_1233, ZN => n_1355);
  g12644 : IND3D0BWP7T port map(A1 => new_item_set, B1 => n_1211, B2 => n_1333, ZN => n_1585);
  g12647 : INVD4BWP7T port map(I => n_1354, ZN => head(3));
  g12649 : INVD4BWP7T port map(I => n_1352, ZN => head(5));
  g12651 : INVD4BWP7T port map(I => n_1351, ZN => head(4));
  g12653 : INVD4BWP7T port map(I => n_1350, ZN => head(0));
  g12655 : INVD4BWP7T port map(I => n_1349, ZN => head(11));
  g12657 : INVD4BWP7T port map(I => n_1348, ZN => head(8));
  g12660 : INVD4BWP7T port map(I => n_1347, ZN => head(2));
  g12662 : INVD4BWP7T port map(I => n_1346, ZN => head(1));
  g12664 : INVD4BWP7T port map(I => n_1345, ZN => head(10));
  g12666 : INVD4BWP7T port map(I => n_1344, ZN => head(9));
  g12668 : INVD4BWP7T port map(I => n_1343, ZN => head(7));
  g12669 : MOAI22D0BWP7T port map(A1 => n_1277, A2 => n_1209, B1 => n_1278, B2 => new_corner(0), ZN => n_1341);
  g12670 : ND2D4BWP7T port map(A1 => n_1304, A2 => n_1279, ZN => clear_tail_flag);
  g12671 : INR4D0BWP7T port map(A1 => n_1740, B1 => corner_count(29), B2 => corner_count(31), B3 => corner_count(30), ZN => n_1340);
  g12672 : OR4D0BWP7T port map(A1 => n_1581, A2 => n_1582, A3 => n_1583, A4 => n_1584, Z => n_1339);
  g12673 : ND4D0BWP7T port map(A1 => n_1286, A2 => n_1252, A3 => n_1240, A4 => n_1250, ZN => n_1338);
  g12675 : INVD4BWP7T port map(I => n_1337, ZN => head(6));
  g12676 : OAI21D0BWP7T port map(A1 => n_1280, A2 => n_1266, B => n_1225, ZN => n_1336);
  g12677 : AO22D0BWP7T port map(A1 => n_1278, A2 => new_corner(5), B1 => new_tail(5), B2 => n_1670, Z => n_1335);
  g12678 : NR2D0BWP7T port map(A1 => n_1307, A2 => send_corner_flag, ZN => n_1334);
  g12679 : AOI21D0BWP7T port map(A1 => n_1570, A2 => n_1217, B => n_1568, ZN => n_1342);
  g12680 : IND3D0BWP7T port map(A1 => n_1718, B1 => n_1276, B2 => n_1282, ZN => n_1386);
  g12681 : AOI211D0BWP7T port map(A1 => n_1264, A2 => n_1578, B => n_1705, C => n_1739, ZN => n_1384);
  g12683 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(7), Z => n_1332);
  g12684 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(0), Z => n_1331);
  g12685 : INR2D0BWP7T port map(A1 => new_item(11), B1 => n_1282, ZN => n_1330);
  g12686 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(1), Z => n_1329);
  g12687 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(2), Z => n_1328);
  g12688 : INR2D0BWP7T port map(A1 => new_item(10), B1 => n_1282, ZN => n_1327);
  g12689 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(4), Z => n_1326);
  g12690 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(5), Z => n_1325);
  g12691 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(6), Z => n_1324);
  g12692 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(8), Z => n_1323);
  g12693 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(9), Z => n_1322);
  g12694 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(10), Z => n_1321);
  g12695 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(11), Z => n_1320);
  g12696 : INR2D0BWP7T port map(A1 => new_item(2), B1 => n_1282, ZN => n_1319);
  g12698 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(3), Z => n_1318);
  g12699 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(9), Z => n_1317);
  g12700 : INR2D0BWP7T port map(A1 => new_item(6), B1 => n_1282, ZN => n_1316);
  g12701 : IND2D0BWP7T port map(A1 => new_head(5), B1 => n_1731, ZN => n_1315);
  g12702 : INR2D0BWP7T port map(A1 => n_1736, B1 => n_1211, ZN => n_1564);
  g12703 : INR2D0BWP7T port map(A1 => n_1662, B1 => n_1211, ZN => n_1565);
  g12704 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(6), Z => n_1314);
  g12705 : IND2D0BWP7T port map(A1 => new_head(4), B1 => n_1731, ZN => n_1313);
  g12706 : IND2D0BWP7T port map(A1 => new_head(0), B1 => n_1731, ZN => n_1312);
  g12707 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(1), Z => n_1311);
  g12708 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(2), Z => n_1310);
  g12709 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(3), Z => n_1309);
  g12710 : AN2D1BWP7T port map(A1 => n_1273, A2 => new_item_set, Z => n_1574);
  g12711 : INR2D0BWP7T port map(A1 => n_1273, B1 => remove_item_set, ZN => n_1333);
  g12712 : CKND1BWP7T port map(I => n_1307, ZN => n_1306);
  g12713 : INVD1BWP7T port map(I => n_1305, ZN => n_1304);
  g12714 : INR2D0BWP7T port map(A1 => new_item(9), B1 => n_1282, ZN => n_1302);
  g12715 : INR2D0BWP7T port map(A1 => new_item(0), B1 => n_1282, ZN => n_1301);
  g12716 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(10), Z => n_1300);
  g12717 : INR2D0BWP7T port map(A1 => new_item(1), B1 => n_1282, ZN => n_1299);
  g12718 : INR2D0BWP7T port map(A1 => new_item(3), B1 => n_1282, ZN => n_1298);
  g12719 : INR2D0BWP7T port map(A1 => new_item(4), B1 => n_1282, ZN => n_1297);
  g12720 : INR2D0BWP7T port map(A1 => new_item(5), B1 => n_1282, ZN => n_1296);
  g12721 : INR2D0BWP7T port map(A1 => new_item(7), B1 => n_1282, ZN => n_1295);
  g12722 : INR2D0BWP7T port map(A1 => new_item(8), B1 => n_1282, ZN => n_1294);
  g12723 : IND2D0BWP7T port map(A1 => new_head(11), B1 => n_1731, ZN => n_1293);
  g12724 : IND2D0BWP7T port map(A1 => new_head(8), B1 => n_1731, ZN => n_1292);
  g12725 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(7), Z => n_1291);
  g12726 : NR4D0BWP7T port map(A1 => n_1247, A2 => n_1248, A3 => n_1261, A4 => n_1251, ZN => n_1290);
  g12727 : ND4D0BWP7T port map(A1 => n_1231, A2 => n_1239, A3 => n_1258, A4 => n_1260, ZN => n_1289);
  g12728 : NR4D0BWP7T port map(A1 => n_1230, A2 => n_1232, A3 => n_1229, A4 => n_1257, ZN => n_1288);
  g12729 : OAI21D0BWP7T port map(A1 => n_1263, A2 => n_1264, B => n_1224, ZN => n_1287);
  g12730 : AOI211D0BWP7T port map(A1 => n_1207, A2 => N(4), B => n_1243, C => n_1259, ZN => n_1286);
  g12731 : ND4D0BWP7T port map(A1 => n_1235, A2 => n_1237, A3 => n_1242, A4 => n_1245, ZN => n_1285);
  g12732 : ND4D0BWP7T port map(A1 => n_1228, A2 => n_1241, A3 => n_1238, A4 => n_1236, ZN => n_1284);
  g12733 : AN4D1BWP7T port map(A1 => n_1255, A2 => n_1253, A3 => n_1254, A4 => n_1256, Z => n_1580);
  g12735 : OR2D0BWP7T port map(A1 => n_1732, A2 => n_1733, Z => n_1579);
  g12736 : ND2D0BWP7T port map(A1 => n_1280, A2 => n_1224, ZN => n_1307);
  g12737 : AOI21D0BWP7T port map(A1 => n_1267, A2 => n_1203, B => n_1216, ZN => n_1305);
  g12738 : OR2D0BWP7T port map(A1 => n_1704, A2 => n_1657, Z => n_1303);
  g12739 : OA21D0BWP7T port map(A1 => n_1263, A2 => n_1265, B => n_1225, Z => n_1569);
  g12740 : OR2D0BWP7T port map(A1 => n_1731, A2 => n_1278, Z => n_1568);
  g12741 : OAI221D0BWP7T port map(A1 => n_1227, A2 => n_1204, B1 => state(1), B2 => state(2), C => n_1224, ZN => n_1651);
  g12742 : ND2D0BWP7T port map(A1 => n_1281, A2 => n_1276, ZN => n_1353);
  g12743 : INVD1BWP7T port map(I => n_1283, ZN => n_1572);
  g12744 : INVD1BWP7T port map(I => n_1281, ZN => n_1731);
  g12745 : AN2D4BWP7T port map(A1 => n_1270, A2 => n_1578, Z => clear_head_flag);
  g12746 : AN2D1BWP7T port map(A1 => n_1265, A2 => n_1225, Z => n_1738);
  g12747 : INR2D0BWP7T port map(A1 => n_1264, B1 => n_1216, ZN => n_1663);
  g12748 : AN2D1BWP7T port map(A1 => n_1264, A2 => n_1224, Z => n_1653);
  g12749 : AN2D1BWP7T port map(A1 => n_1202, A2 => n_1273, Z => n_1575);
  g12750 : OR2D0BWP7T port map(A1 => n_1266, A2 => n_1264, Z => n_1570);
  g12751 : NR2XD0BWP7T port map(A1 => n_1203, A2 => n_1216, ZN => n_1703);
  g12752 : NR2D0BWP7T port map(A1 => n_1269, A2 => n_1226, ZN => n_1734);
  g12753 : AN2D1BWP7T port map(A1 => n_1266, A2 => n_1224, Z => n_1732);
  g12754 : INR2D0BWP7T port map(A1 => n_1266, B1 => n_1216, ZN => n_1654);
  g12756 : NR2D0BWP7T port map(A1 => n_1272, A2 => n_1216, ZN => n_1657);
  g12757 : AN2D1BWP7T port map(A1 => n_1264, A2 => n_1225, Z => n_1733);
  g12758 : ND2D0BWP7T port map(A1 => n_1265, A2 => n_1217, ZN => n_1283);
  g12759 : ND2D0BWP7T port map(A1 => n_1266, A2 => n_1578, ZN => n_1282);
  g12760 : ND2D0BWP7T port map(A1 => n_1263, A2 => n_1217, ZN => n_1281);
  g12761 : CKND1BWP7T port map(I => n_1670, ZN => n_1277);
  g12762 : INVD0BWP7T port map(I => n_1739, ZN => n_1276);
  g12763 : INR2D0BWP7T port map(A1 => n_1263, B1 => n_1226, ZN => n_1735);
  g12764 : OAI211D0BWP7T port map(A1 => state(3), A2 => n_1205, B => state(2), C => state(4), ZN => n_1275);
  g12765 : NR4D0BWP7T port map(A1 => new_tail(4), A2 => new_tail(3), A3 => new_tail(2), A4 => new_tail(1), ZN => n_1274);
  g12766 : NR2D0BWP7T port map(A1 => n_1267, A2 => n_1223, ZN => n_1662);
  g12767 : INR2D0BWP7T port map(A1 => n_1263, B1 => n_1222, ZN => n_1718);
  g12768 : ND2D0BWP7T port map(A1 => n_1267, A2 => n_1272, ZN => n_1280);
  g12769 : AN2D2BWP7T port map(A1 => n_1268, A2 => n_1578, Z => n_1704);
  g12770 : NR2D0BWP7T port map(A1 => n_1272, A2 => n_1223, ZN => n_1736);
  g12771 : OR4D0BWP7T port map(A1 => n_146, A2 => n_1701, A3 => n_1700, A4 => n_1699, Z => n_1581);
  g12772 : AN2D4BWP7T port map(A1 => n_1271, A2 => n_1578, Z => clear_corner_flag);
  g12773 : AN2D1BWP7T port map(A1 => n_1263, A2 => n_1224, Z => n_1737);
  g12774 : AN2D4BWP7T port map(A1 => n_1268, A2 => n_1224, Z => new_item_clear);
  g12775 : ND2D1BWP7T port map(A1 => n_1265, A2 => n_1224, ZN => n_1279);
  g12776 : INR2D0BWP7T port map(A1 => n_1265, B1 => n_1222, ZN => n_1278);
  g12777 : NR2XD0BWP7T port map(A1 => n_1267, A2 => n_1216, ZN => n_1670);
  g12778 : NR2XD0BWP7T port map(A1 => n_1269, A2 => n_1216, ZN => n_1739);
  g12779 : NR2D0BWP7T port map(A1 => n_1267, A2 => n_1222, ZN => n_1705);
  g12780 : INVD0BWP7T port map(I => n_1271, ZN => n_1272);
  g12781 : INVD0BWP7T port map(I => n_1203, ZN => n_1270);
  g12782 : INVD1BWP7T port map(I => n_1269, ZN => n_1268);
  g12783 : MAOI22D0BWP7T port map(A1 => n_1214, A2 => N(5), B1 => n_1207, B2 => N(4), ZN => n_1262);
  g12784 : CKXOR2D0BWP7T port map(A1 => N(14), A2 => corner_count(14), Z => n_1261);
  g12785 : XNR2D1BWP7T port map(A1 => corner_count(8), A2 => N(8), ZN => n_1260);
  g12786 : CKXOR2D0BWP7T port map(A1 => N(29), A2 => corner_count(29), Z => n_1259);
  g12787 : XNR2D1BWP7T port map(A1 => corner_count(9), A2 => N(9), ZN => n_1258);
  g12788 : CKXOR2D0BWP7T port map(A1 => N(16), A2 => corner_count(16), Z => n_1257);
  g12789 : NR4D0BWP7T port map(A1 => n_1683, A2 => n_1684, A3 => n_1685, A4 => n_1686, ZN => n_1256);
  g12790 : NR4D0BWP7T port map(A1 => n_1671, A2 => n_1672, A3 => n_1673, A4 => n_1674, ZN => n_1255);
  g12791 : NR4D0BWP7T port map(A1 => n_1679, A2 => n_1680, A3 => n_1681, A4 => n_1682, ZN => n_1254);
  g12792 : NR4D0BWP7T port map(A1 => n_1675, A2 => n_1676, A3 => n_1677, A4 => n_1678, ZN => n_1253);
  g12793 : INR3D0BWP7T port map(A1 => remove_item_set, B1 => remove_item_type, B2 => new_item_set, ZN => n_1742);
  g12794 : AOI22D0BWP7T port map(A1 => corner_count(5), A2 => n_1208, B1 => n_1206, B2 => N(6), ZN => n_1252);
  g12795 : OR4D0BWP7T port map(A1 => n_1690, A2 => n_1689, A3 => n_1688, A4 => n_1687, Z => n_1584);
  g12796 : OR4D0BWP7T port map(A1 => n_1694, A2 => n_1693, A3 => n_1692, A4 => n_1691, Z => n_1583);
  g12797 : OR4D0BWP7T port map(A1 => n_1698, A2 => n_1697, A3 => n_1696, A4 => n_1695, Z => n_1582);
  g12799 : NR3D0BWP7T port map(A1 => new_head_flag, A2 => new_corner_flag, A3 => new_tail_flag, ZN => n_1273);
  g12800 : NR2XD0BWP7T port map(A1 => n_1221, A2 => n_1204, ZN => n_1271);
  g12802 : ND2D1BWP7T port map(A1 => n_1227, A2 => n_1204, ZN => n_1269);
  g12803 : ND2D1BWP7T port map(A1 => n_1218, A2 => state(2), ZN => n_1267);
  g12804 : INR2D0BWP7T port map(A1 => n_1227, B1 => n_1204, ZN => n_1266);
  g12805 : NR2XD0BWP7T port map(A1 => n_1219, A2 => state(2), ZN => n_1265);
  g12806 : NR2D0BWP7T port map(A1 => n_1221, A2 => state(2), ZN => n_1264);
  g12807 : NR2D0BWP7T port map(A1 => n_1220, A2 => state(2), ZN => n_1263);
  g12808 : CKXOR2D0BWP7T port map(A1 => N(12), A2 => corner_count(12), Z => n_1251);
  g12809 : XNR2D1BWP7T port map(A1 => corner_count(28), A2 => N(28), ZN => n_1250);
  g12810 : CKXOR2D0BWP7T port map(A1 => N(7), A2 => corner_count(7), Z => n_1249);
  g12811 : CKXOR2D0BWP7T port map(A1 => N(15), A2 => corner_count(15), Z => n_1248);
  g12812 : CKXOR2D0BWP7T port map(A1 => N(13), A2 => corner_count(13), Z => n_1247);
  g12813 : CKXOR2D0BWP7T port map(A1 => N(27), A2 => corner_count(27), Z => n_1246);
  g12814 : XNR2D1BWP7T port map(A1 => corner_count(3), A2 => N(3), ZN => n_1245);
  g12815 : CKXOR2D0BWP7T port map(A1 => N(25), A2 => corner_count(25), Z => n_1244);
  g12816 : CKXOR2D0BWP7T port map(A1 => N(31), A2 => corner_count(31), Z => n_1243);
  g12817 : XNR2D1BWP7T port map(A1 => corner_count(2), A2 => N(2), ZN => n_1242);
  g12818 : XNR2D1BWP7T port map(A1 => corner_count(21), A2 => N(21), ZN => n_1241);
  g12819 : XNR2D1BWP7T port map(A1 => corner_count(30), A2 => N(30), ZN => n_1240);
  g12820 : XNR2D1BWP7T port map(A1 => corner_count(10), A2 => N(10), ZN => n_1239);
  g12821 : XNR2D1BWP7T port map(A1 => corner_count(23), A2 => N(23), ZN => n_1238);
  g12822 : MAOI22D0BWP7T port map(A1 => n_1212, A2 => N(1), B1 => n_1212, B2 => N(1), ZN => n_1237);
  g12823 : XNR2D1BWP7T port map(A1 => corner_count(20), A2 => N(20), ZN => n_1236);
  g12824 : AOI22D0BWP7T port map(A1 => corner_count(0), A2 => n_152, B1 => n_146, B2 => N(0), ZN => n_1235);
  g12825 : XNR2D1BWP7T port map(A1 => corner_count(26), A2 => N(26), ZN => n_1234);
  g12826 : XNR2D1BWP7T port map(A1 => corner_count(24), A2 => N(24), ZN => n_1233);
  g12827 : CKXOR2D0BWP7T port map(A1 => N(19), A2 => corner_count(19), Z => n_1232);
  g12828 : XNR2D1BWP7T port map(A1 => corner_count(11), A2 => N(11), ZN => n_1231);
  g12829 : CKXOR2D0BWP7T port map(A1 => N(18), A2 => corner_count(18), Z => n_1230);
  g12830 : CKXOR2D0BWP7T port map(A1 => N(17), A2 => corner_count(17), Z => n_1229);
  g12831 : XNR2D1BWP7T port map(A1 => corner_count(22), A2 => N(22), ZN => n_1228);
  g12832 : MOAI22D0BWP7T port map(A1 => corner_count(1), A2 => corner_count(2), B1 => corner_count(1), B2 => corner_count(2), ZN => n_1740);
  g12833 : INVD0BWP7T port map(I => n_1226, ZN => n_1225);
  g12834 : INVD0BWP7T port map(I => n_1224, ZN => n_1223);
  g12835 : INVD0BWP7T port map(I => n_1578, ZN => n_1222);
  g12836 : NR2XD0BWP7T port map(A1 => state(0), A2 => state(1), ZN => n_1227);
  g12837 : ND2D0BWP7T port map(A1 => state(3), A2 => state(4), ZN => n_1226);
  g12838 : INR2XD0BWP7T port map(A1 => state(4), B1 => state(3), ZN => n_1224);
  g12839 : INR2XD0BWP7T port map(A1 => state(3), B1 => state(4), ZN => n_1578);
  g12841 : INVD0BWP7T port map(I => n_1218, ZN => n_1219);
  g12842 : INVD1BWP7T port map(I => n_1217, ZN => n_1216);
  g12843 : IND2D0BWP7T port map(A1 => N(6), B1 => corner_count(6), ZN => n_1215);
  g12844 : ND2D1BWP7T port map(A1 => state(1), A2 => state(0), ZN => n_1221);
  g12845 : ND2D1BWP7T port map(A1 => n_1205, A2 => state(1), ZN => n_1220);
  g12846 : NR2XD0BWP7T port map(A1 => n_1205, A2 => state(1), ZN => n_1218);
  g12847 : NR2XD0BWP7T port map(A1 => state(4), A2 => state(3), ZN => n_1217);
  g12848 : CKND1BWP7T port map(I => corner_count(5), ZN => n_1214);
  g12850 : INVD0BWP7T port map(I => corner_count(1), ZN => n_1212);
  g12853 : INVD1BWP7T port map(I => send_corner_flag, ZN => n_1211);
  g12854 : INVD0BWP7T port map(I => new_head_flag, ZN => n_1210);
  g12855 : CKND1BWP7T port map(I => new_tail(0), ZN => n_1209);
  g12856 : CKND1BWP7T port map(I => N(5), ZN => n_1208);
  g12857 : CKND1BWP7T port map(I => corner_count(4), ZN => n_1207);
  g12858 : CKND1BWP7T port map(I => corner_count(6), ZN => n_1206);
  g2 : INR3D0BWP7T port map(A1 => n_1333, B1 => new_item_set, B2 => n_1211, ZN => n_1573);
  g12861 : IND2D1BWP7T port map(A1 => n_1220, B1 => state(2), ZN => n_1203);
  g12862 : INR3D0BWP7T port map(A1 => new_item_set, B1 => new_item(0), B2 => new_item(1), ZN => n_1202);
  N_reg_0 : LNQD1BWP7T port map(EN => n_483, D => n_190, Q => N(0));
  N_reg_1 : LNQD1BWP7T port map(EN => n_483, D => n_162, Q => N(1));
  N_reg_2 : LNQD1BWP7T port map(EN => n_483, D => n_163, Q => N(2));
  N_reg_3 : LNQD1BWP7T port map(EN => n_483, D => n_191, Q => N(3));
  N_reg_4 : LNQD1BWP7T port map(EN => n_483, D => n_165, Q => N(4));
  N_reg_5 : LNQD1BWP7T port map(EN => n_483, D => n_169, Q => N(5));
  N_reg_6 : LNQD1BWP7T port map(EN => n_483, D => n_170, Q => N(6));
  N_reg_7 : LNQD1BWP7T port map(EN => n_483, D => n_173, Q => N(7));
  N_reg_8 : LNQD1BWP7T port map(EN => n_483, D => n_160, Q => N(8));
  N_reg_9 : LNQD1BWP7T port map(EN => n_483, D => n_159, Q => N(9));
  N_reg_10 : LNQD1BWP7T port map(EN => n_483, D => n_174, Q => N(10));
  N_reg_11 : LNQD1BWP7T port map(EN => n_483, D => n_167, Q => N(11));
  N_reg_12 : LNQD1BWP7T port map(EN => n_483, D => n_172, Q => N(12));
  N_reg_13 : LNQD1BWP7T port map(EN => n_483, D => n_178, Q => N(13));
  N_reg_14 : LNQD1BWP7T port map(EN => n_483, D => n_175, Q => N(14));
  N_reg_15 : LNQD1BWP7T port map(EN => n_483, D => n_177, Q => N(15));
  N_reg_16 : LNQD1BWP7T port map(EN => n_483, D => n_180, Q => N(16));
  N_reg_17 : LNQD1BWP7T port map(EN => n_483, D => n_166, Q => N(17));
  N_reg_18 : LNQD1BWP7T port map(EN => n_483, D => n_176, Q => N(18));
  N_reg_19 : LNQD1BWP7T port map(EN => n_483, D => n_179, Q => N(19));
  N_reg_20 : LNQD1BWP7T port map(EN => n_483, D => n_181, Q => N(20));
  N_reg_21 : LNQD1BWP7T port map(EN => n_483, D => n_171, Q => N(21));
  N_reg_22 : LNQD1BWP7T port map(EN => n_483, D => n_161, Q => N(22));
  N_reg_23 : LNQD1BWP7T port map(EN => n_483, D => n_158, Q => N(23));
  N_reg_24 : LNQD1BWP7T port map(EN => n_483, D => n_183, Q => N(24));
  N_reg_25 : LNQD1BWP7T port map(EN => n_483, D => n_168, Q => N(25));
  N_reg_26 : LNQD1BWP7T port map(EN => n_483, D => n_184, Q => N(26));
  N_reg_27 : LNQD1BWP7T port map(EN => n_483, D => n_185, Q => N(27));
  N_reg_28 : LNQD1BWP7T port map(EN => n_483, D => n_186, Q => N(28));
  N_reg_29 : LNQD1BWP7T port map(EN => n_483, D => n_182, Q => N(29));
  N_reg_30 : LNQD1BWP7T port map(EN => n_483, D => n_188, Q => N(30));
  N_reg_31 : LNQD1BWP7T port map(EN => n_483, D => n_189, Q => N(31));
  S_S_reg_1_0 : LHQD1BWP7T port map(E => n_674, D => n_279, Q => n_1180);
  S_S_reg_1_1 : LHQD1BWP7T port map(E => n_674, D => n_393, Q => n_1181);
  S_S_reg_1_2 : LHQD1BWP7T port map(E => n_674, D => n_388, Q => n_1182);
  S_S_reg_1_3 : LHQD1BWP7T port map(E => n_674, D => n_386, Q => n_1183);
  S_S_reg_1_4 : LHQD1BWP7T port map(E => n_674, D => n_381, Q => n_1184);
  S_S_reg_1_5 : LHQD1BWP7T port map(E => n_674, D => n_374, Q => n_1185);
  S_S_reg_2_0 : LHQD1BWP7T port map(E => n_764, D => n_376, Q => n_1174);
  S_S_reg_2_1 : LHQD1BWP7T port map(E => n_764, D => n_348, Q => n_1175);
  S_S_reg_2_2 : LHQD1BWP7T port map(E => n_764, D => n_370, Q => n_1176);
  S_S_reg_2_3 : LHQD1BWP7T port map(E => n_764, D => n_367, Q => n_1177);
  S_S_reg_2_4 : LHQD1BWP7T port map(E => n_764, D => n_363, Q => n_1178);
  S_S_reg_2_5 : LHQD1BWP7T port map(E => n_764, D => n_410, Q => n_1179);
  S_S_reg_3_0 : LHQD1BWP7T port map(E => n_766, D => n_396, Q => n_1168);
  S_S_reg_3_1 : LHQD1BWP7T port map(E => n_766, D => n_353, Q => n_1169);
  S_S_reg_3_2 : LHQD1BWP7T port map(E => n_766, D => n_355, Q => n_1170);
  S_S_reg_3_3 : LHQD1BWP7T port map(E => n_766, D => n_294, Q => n_1171);
  S_S_reg_3_4 : LHQD1BWP7T port map(E => n_766, D => n_352, Q => n_1172);
  S_S_reg_3_5 : LHQD1BWP7T port map(E => n_766, D => n_350, Q => n_1173);
  S_S_reg_4_0 : LNQD1BWP7T port map(EN => n_598, D => n_349, Q => n_1162);
  S_S_reg_4_1 : LNQD1BWP7T port map(EN => n_598, D => n_298, Q => n_1163);
  S_S_reg_4_2 : LNQD1BWP7T port map(EN => n_598, D => n_345, Q => n_1164);
  S_S_reg_4_3 : LNQD1BWP7T port map(EN => n_598, D => n_344, Q => n_1165);
  S_S_reg_4_4 : LNQD1BWP7T port map(EN => n_598, D => n_343, Q => n_1166);
  S_S_reg_4_5 : LNQD1BWP7T port map(EN => n_598, D => n_356, Q => n_1167);
  S_S_reg_5_0 : LNQD1BWP7T port map(EN => n_673, D => n_394, Q => n_1156);
  S_S_reg_5_1 : LNQD1BWP7T port map(EN => n_673, D => n_401, Q => n_1157);
  S_S_reg_5_2 : LNQD1BWP7T port map(EN => n_673, D => n_398, Q => n_1158);
  S_S_reg_5_3 : LNQD1BWP7T port map(EN => n_673, D => n_335, Q => n_1159);
  S_S_reg_5_4 : LNQD1BWP7T port map(EN => n_673, D => n_395, Q => n_1160);
  S_S_reg_5_5 : LNQD1BWP7T port map(EN => n_673, D => n_375, Q => n_1161);
  S_S_reg_6_0 : LHQD1BWP7T port map(E => n_765, D => n_321, Q => n_1150);
  S_S_reg_6_1 : LHQD1BWP7T port map(E => n_765, D => n_284, Q => n_1151);
  S_S_reg_6_2 : LHQD1BWP7T port map(E => n_765, D => n_286, Q => n_1152);
  S_S_reg_6_3 : LHQD1BWP7T port map(E => n_765, D => n_413, Q => n_1153);
  S_S_reg_6_4 : LHQD1BWP7T port map(E => n_765, D => n_354, Q => n_1154);
  S_S_reg_6_5 : LHQD1BWP7T port map(E => n_765, D => n_288, Q => n_1155);
  S_S_reg_7_0 : LHQD1BWP7T port map(E => n_763, D => n_406, Q => n_1144);
  S_S_reg_7_1 : LHQD1BWP7T port map(E => n_763, D => n_399, Q => n_1145);
  S_S_reg_7_2 : LHQD1BWP7T port map(E => n_763, D => n_402, Q => n_1146);
  S_S_reg_7_3 : LHQD1BWP7T port map(E => n_763, D => n_403, Q => n_1147);
  S_S_reg_7_4 : LHQD1BWP7T port map(E => n_763, D => n_404, Q => n_1148);
  S_S_reg_7_5 : LHQD1BWP7T port map(E => n_763, D => n_308, Q => n_1149);
  S_S_reg_8_0 : LNQD1BWP7T port map(EN => n_762, D => n_342, Q => n_1138);
  S_S_reg_8_1 : LNQD1BWP7T port map(EN => n_762, D => n_405, Q => n_1139);
  S_S_reg_8_2 : LNQD1BWP7T port map(EN => n_762, D => n_319, Q => n_1140);
  S_S_reg_8_3 : LNQD1BWP7T port map(EN => n_762, D => n_408, Q => n_1141);
  S_S_reg_8_4 : LNQD1BWP7T port map(EN => n_762, D => n_409, Q => n_1142);
  S_S_reg_8_5 : LNQD1BWP7T port map(EN => n_762, D => n_411, Q => n_1143);
  S_S_reg_9_0 : LNQD1BWP7T port map(EN => n_761, D => n_397, Q => n_1132);
  S_S_reg_9_1 : LNQD1BWP7T port map(EN => n_761, D => n_412, Q => n_1133);
  S_S_reg_9_2 : LNQD1BWP7T port map(EN => n_761, D => n_400, Q => n_1134);
  S_S_reg_9_3 : LNQD1BWP7T port map(EN => n_761, D => n_414, Q => n_1135);
  S_S_reg_9_4 : LNQD1BWP7T port map(EN => n_761, D => n_360, Q => n_1136);
  S_S_reg_9_5 : LNQD1BWP7T port map(EN => n_761, D => n_415, Q => n_1137);
  S_S_reg_10_0 : LNQD1BWP7T port map(EN => n_760, D => n_328, Q => n_1126);
  S_S_reg_10_1 : LNQD1BWP7T port map(EN => n_760, D => n_416, Q => n_1127);
  S_S_reg_10_2 : LNQD1BWP7T port map(EN => n_760, D => n_340, Q => n_1128);
  S_S_reg_10_3 : LNQD1BWP7T port map(EN => n_760, D => n_339, Q => n_1129);
  S_S_reg_10_4 : LNQD1BWP7T port map(EN => n_760, D => n_338, Q => n_1130);
  S_S_reg_10_5 : LNQD1BWP7T port map(EN => n_760, D => n_337, Q => n_1131);
  S_S_reg_11_0 : LNQD1BWP7T port map(EN => n_759, D => n_336, Q => n_1120);
  S_S_reg_11_1 : LNQD1BWP7T port map(EN => n_759, D => n_334, Q => n_1121);
  S_S_reg_11_2 : LNQD1BWP7T port map(EN => n_759, D => n_333, Q => n_1122);
  S_S_reg_11_3 : LNQD1BWP7T port map(EN => n_759, D => n_332, Q => n_1123);
  S_S_reg_11_4 : LNQD1BWP7T port map(EN => n_759, D => n_331, Q => n_1124);
  S_S_reg_11_5 : LNQD1BWP7T port map(EN => n_759, D => n_330, Q => n_1125);
  S_S_reg_12_0 : LNQD1BWP7T port map(EN => n_758, D => n_329, Q => n_1114);
  S_S_reg_12_1 : LNQD1BWP7T port map(EN => n_758, D => n_327, Q => n_1115);
  S_S_reg_12_2 : LNQD1BWP7T port map(EN => n_758, D => n_326, Q => n_1116);
  S_S_reg_12_3 : LNQD1BWP7T port map(EN => n_758, D => n_325, Q => n_1117);
  S_S_reg_12_4 : LNQD1BWP7T port map(EN => n_758, D => n_324, Q => n_1118);
  S_S_reg_12_5 : LNQD1BWP7T port map(EN => n_758, D => n_323, Q => n_1119);
  S_S_reg_13_0 : LNQD1BWP7T port map(EN => n_757, D => n_322, Q => n_1108);
  S_S_reg_13_1 : LNQD1BWP7T port map(EN => n_757, D => n_320, Q => n_1109);
  S_S_reg_13_2 : LNQD1BWP7T port map(EN => n_757, D => n_318, Q => n_1110);
  S_S_reg_13_3 : LNQD1BWP7T port map(EN => n_757, D => n_317, Q => n_1111);
  S_S_reg_13_4 : LNQD1BWP7T port map(EN => n_757, D => n_316, Q => n_1112);
  S_S_reg_13_5 : LNQD1BWP7T port map(EN => n_757, D => n_315, Q => n_1113);
  S_S_reg_14_0 : LHQD1BWP7T port map(E => n_756, D => n_314, Q => n_1102);
  S_S_reg_14_1 : LHQD1BWP7T port map(E => n_756, D => n_313, Q => n_1103);
  S_S_reg_14_2 : LHQD1BWP7T port map(E => n_756, D => n_312, Q => n_1104);
  S_S_reg_14_3 : LHQD1BWP7T port map(E => n_756, D => n_311, Q => n_1105);
  S_S_reg_14_4 : LHQD1BWP7T port map(E => n_756, D => n_310, Q => n_1106);
  S_S_reg_14_5 : LHQD1BWP7T port map(E => n_756, D => n_309, Q => n_1107);
  S_S_reg_15_0 : LHQD1BWP7T port map(E => n_702, D => n_307, Q => n_1096);
  S_S_reg_15_1 : LHQD1BWP7T port map(E => n_702, D => n_306, Q => n_1097);
  S_S_reg_15_2 : LHQD1BWP7T port map(E => n_702, D => n_305, Q => n_1098);
  S_S_reg_15_3 : LHQD1BWP7T port map(E => n_702, D => n_304, Q => n_1099);
  S_S_reg_15_4 : LHQD1BWP7T port map(E => n_702, D => n_303, Q => n_1100);
  S_S_reg_15_5 : LHQD1BWP7T port map(E => n_702, D => n_302, Q => n_1101);
  S_S_reg_16_0 : LHQD1BWP7T port map(E => n_812, D => n_301, Q => n_1090);
  S_S_reg_16_1 : LHQD1BWP7T port map(E => n_812, D => n_300, Q => n_1091);
  S_S_reg_16_2 : LHQD1BWP7T port map(E => n_812, D => n_299, Q => n_1092);
  S_S_reg_16_3 : LHQD1BWP7T port map(E => n_812, D => n_297, Q => n_1093);
  S_S_reg_16_4 : LHQD1BWP7T port map(E => n_812, D => n_296, Q => n_1094);
  S_S_reg_16_5 : LHQD1BWP7T port map(E => n_812, D => n_295, Q => n_1095);
  S_S_reg_17_0 : LHQD1BWP7T port map(E => n_859, D => n_407, Q => n_1084);
  S_S_reg_17_1 : LHQD1BWP7T port map(E => n_859, D => n_293, Q => n_1085);
  S_S_reg_17_2 : LHQD1BWP7T port map(E => n_859, D => n_292, Q => n_1086);
  S_S_reg_17_3 : LHQD1BWP7T port map(E => n_859, D => n_291, Q => n_1087);
  S_S_reg_17_4 : LHQD1BWP7T port map(E => n_859, D => n_290, Q => n_1088);
  S_S_reg_17_5 : LHQD1BWP7T port map(E => n_859, D => n_289, Q => n_1089);
  S_S_reg_18_0 : LNQD1BWP7T port map(EN => n_887, D => n_287, Q => n_1078);
  S_S_reg_18_1 : LNQD1BWP7T port map(EN => n_887, D => n_285, Q => n_1079);
  S_S_reg_18_2 : LNQD1BWP7T port map(EN => n_887, D => n_283, Q => n_1080);
  S_S_reg_18_3 : LNQD1BWP7T port map(EN => n_887, D => n_282, Q => n_1081);
  S_S_reg_18_4 : LNQD1BWP7T port map(EN => n_887, D => n_281, Q => n_1082);
  S_S_reg_18_5 : LNQD1BWP7T port map(EN => n_887, D => n_280, Q => n_1083);
  S_S_reg_19_0 : LNQD1BWP7T port map(EN => n_886, D => n_278, Q => n_1072);
  S_S_reg_19_1 : LNQD1BWP7T port map(EN => n_886, D => n_277, Q => n_1073);
  S_S_reg_19_2 : LNQD1BWP7T port map(EN => n_886, D => n_276, Q => n_1074);
  S_S_reg_19_3 : LNQD1BWP7T port map(EN => n_886, D => n_275, Q => n_1075);
  S_S_reg_19_4 : LNQD1BWP7T port map(EN => n_886, D => n_274, Q => n_1076);
  S_S_reg_19_5 : LNQD1BWP7T port map(EN => n_886, D => n_273, Q => n_1077);
  S_S_reg_20_0 : LHQD1BWP7T port map(E => n_811, D => n_392, Q => n_1066);
  S_S_reg_20_1 : LHQD1BWP7T port map(E => n_811, D => n_391, Q => n_1067);
  S_S_reg_20_2 : LHQD1BWP7T port map(E => n_811, D => n_390, Q => n_1068);
  S_S_reg_20_3 : LHQD1BWP7T port map(E => n_811, D => n_389, Q => n_1069);
  S_S_reg_20_4 : LHQD1BWP7T port map(E => n_811, D => n_387, Q => n_1070);
  S_S_reg_20_5 : LHQD1BWP7T port map(E => n_811, D => n_385, Q => n_1071);
  S_S_reg_21_0 : LNQD1BWP7T port map(EN => n_860, D => n_384, Q => n_1060);
  S_S_reg_21_1 : LNQD1BWP7T port map(EN => n_860, D => n_383, Q => n_1061);
  S_S_reg_21_2 : LNQD1BWP7T port map(EN => n_860, D => n_382, Q => n_1062);
  S_S_reg_21_3 : LNQD1BWP7T port map(EN => n_860, D => n_380, Q => n_1063);
  S_S_reg_21_4 : LNQD1BWP7T port map(EN => n_860, D => n_379, Q => n_1064);
  S_S_reg_21_5 : LNQD1BWP7T port map(EN => n_860, D => n_378, Q => n_1065);
  S_S_reg_22_0 : LHQD1BWP7T port map(E => n_889, D => n_377, Q => n_1054);
  S_S_reg_22_1 : LHQD1BWP7T port map(E => n_889, D => n_373, Q => n_1055);
  S_S_reg_22_2 : LHQD1BWP7T port map(E => n_889, D => n_372, Q => n_1056);
  S_S_reg_22_3 : LHQD1BWP7T port map(E => n_889, D => n_371, Q => n_1057);
  S_S_reg_22_4 : LHQD1BWP7T port map(E => n_889, D => n_346, Q => n_1058);
  S_S_reg_22_5 : LHQD1BWP7T port map(E => n_889, D => n_347, Q => n_1059);
  S_S_reg_23_0 : LHQD1BWP7T port map(E => n_888, D => n_369, Q => n_1048);
  S_S_reg_23_1 : LHQD1BWP7T port map(E => n_888, D => n_368, Q => n_1049);
  S_S_reg_23_2 : LHQD1BWP7T port map(E => n_888, D => n_366, Q => n_1050);
  S_S_reg_23_3 : LHQD1BWP7T port map(E => n_888, D => n_341, Q => n_1051);
  S_S_reg_23_4 : LHQD1BWP7T port map(E => n_888, D => n_365, Q => n_1052);
  S_S_reg_23_5 : LHQD1BWP7T port map(E => n_888, D => n_364, Q => n_1053);
  S_S_reg_24_0 : LHQD1BWP7T port map(E => n_890, D => n_362, Q => n_1042);
  S_S_reg_24_1 : LHQD1BWP7T port map(E => n_890, D => n_361, Q => n_1043);
  S_S_reg_24_2 : LHQD1BWP7T port map(E => n_890, D => n_351, Q => n_1044);
  S_S_reg_24_3 : LHQD1BWP7T port map(E => n_890, D => n_358, Q => n_1045);
  S_S_reg_24_4 : LHQD1BWP7T port map(E => n_890, D => n_359, Q => n_1046);
  S_S_reg_24_5 : LHQD1BWP7T port map(E => n_890, D => n_357, Q => n_1047);
  corner_check_reg_5 : LNQD1BWP7T port map(EN => n_530, D => n_1037, Q => corner_check(5));
  corner_count_reg_0 : LNQD1BWP7T port map(EN => n_470, D => n_451, Q => corner_count(0));
  corner_count_reg_1 : LNQD1BWP7T port map(EN => n_470, D => n_251, Q => corner_count(1));
  corner_count_reg_2 : LNQD1BWP7T port map(EN => n_470, D => n_269, Q => corner_count(2));
  corner_count_reg_3 : LNQD1BWP7T port map(EN => n_470, D => n_268, Q => corner_count(3));
  corner_count_reg_4 : LNQD1BWP7T port map(EN => n_470, D => n_270, Q => corner_count(4));
  corner_count_reg_5 : LNQD1BWP7T port map(EN => n_470, D => n_267, Q => corner_count(5));
  corner_count_reg_6 : LNQD1BWP7T port map(EN => n_470, D => n_266, Q => corner_count(6));
  corner_count_reg_7 : LNQD1BWP7T port map(EN => n_470, D => n_265, Q => corner_count(7));
  corner_count_reg_8 : LNQD1BWP7T port map(EN => n_470, D => n_264, Q => corner_count(8));
  corner_count_reg_9 : LNQD1BWP7T port map(EN => n_470, D => n_272, Q => corner_count(9));
  corner_count_reg_10 : LNQD1BWP7T port map(EN => n_470, D => n_271, Q => corner_count(10));
  corner_count_reg_11 : LNQD1BWP7T port map(EN => n_470, D => n_262, Q => corner_count(11));
  corner_count_reg_12 : LNQD1BWP7T port map(EN => n_470, D => n_250, Q => corner_count(12));
  corner_count_reg_13 : LNQD1BWP7T port map(EN => n_470, D => n_261, Q => corner_count(13));
  corner_count_reg_14 : LNQD1BWP7T port map(EN => n_470, D => n_247, Q => corner_count(14));
  corner_count_reg_15 : LNQD1BWP7T port map(EN => n_470, D => n_242, Q => corner_count(15));
  corner_count_reg_16 : LNQD1BWP7T port map(EN => n_470, D => n_241, Q => corner_count(16));
  corner_count_reg_17 : LNQD1BWP7T port map(EN => n_470, D => n_253, Q => corner_count(17));
  corner_count_reg_18 : LNQD1BWP7T port map(EN => n_470, D => n_260, Q => corner_count(18));
  corner_count_reg_19 : LNQD1BWP7T port map(EN => n_470, D => n_259, Q => corner_count(19));
  corner_count_reg_20 : LNQD1BWP7T port map(EN => n_470, D => n_244, Q => corner_count(20));
  corner_count_reg_21 : LNQD1BWP7T port map(EN => n_470, D => n_248, Q => corner_count(21));
  corner_count_reg_22 : LNQD1BWP7T port map(EN => n_470, D => n_263, Q => corner_count(22));
  corner_count_reg_23 : LNQD1BWP7T port map(EN => n_470, D => n_258, Q => corner_count(23));
  corner_count_reg_24 : LNQD1BWP7T port map(EN => n_470, D => n_243, Q => corner_count(24));
  corner_count_reg_25 : LNQD1BWP7T port map(EN => n_470, D => n_245, Q => corner_count(25));
  corner_count_reg_26 : LNQD1BWP7T port map(EN => n_470, D => n_257, Q => corner_count(26));
  corner_count_reg_27 : LNQD1BWP7T port map(EN => n_470, D => n_256, Q => corner_count(27));
  corner_count_reg_28 : LNQD1BWP7T port map(EN => n_470, D => n_246, Q => corner_count(28));
  corner_count_reg_29 : LNQD1BWP7T port map(EN => n_470, D => n_249, Q => corner_count(29));
  corner_count_reg_30 : LNQD1BWP7T port map(EN => n_470, D => n_255, Q => corner_count(30));
  corner_count_reg_31 : LNQD1BWP7T port map(EN => n_470, D => n_252, Q => corner_count(31));
  new_N_reg_1 : LNQD1BWP7T port map(EN => n_1651, D => n_1617, Q => new_N(1));
  new_N_reg_2 : LNQD1BWP7T port map(EN => n_1651, D => n_1616, Q => new_N(2));
  new_N_reg_3 : LNQD1BWP7T port map(EN => n_1651, D => n_1615, Q => new_N(3));
  new_N_reg_4 : LNQD1BWP7T port map(EN => n_1651, D => n_1614, Q => new_N(4));
  new_N_reg_5 : LNQD1BWP7T port map(EN => n_1651, D => n_1613, Q => new_N(5));
  new_N_reg_6 : LNQD1BWP7T port map(EN => n_1651, D => n_1612, Q => new_N(6));
  new_N_reg_7 : LNQD1BWP7T port map(EN => n_1651, D => n_1611, Q => new_N(7));
  new_N_reg_8 : LNQD1BWP7T port map(EN => n_1651, D => n_1610, Q => new_N(8));
  new_N_reg_9 : LNQD1BWP7T port map(EN => n_1651, D => n_1609, Q => new_N(9));
  new_N_reg_10 : LNQD1BWP7T port map(EN => n_1651, D => n_1608, Q => new_N(10));
  new_N_reg_11 : LNQD1BWP7T port map(EN => n_1651, D => n_1607, Q => new_N(11));
  new_N_reg_12 : LNQD1BWP7T port map(EN => n_1651, D => n_1606, Q => new_N(12));
  new_N_reg_13 : LNQD1BWP7T port map(EN => n_1651, D => n_1605, Q => new_N(13));
  new_N_reg_14 : LNQD1BWP7T port map(EN => n_1651, D => n_1604, Q => new_N(14));
  new_N_reg_15 : LNQD1BWP7T port map(EN => n_1651, D => n_1603, Q => new_N(15));
  new_N_reg_16 : LNQD1BWP7T port map(EN => n_1651, D => n_1602, Q => new_N(16));
  new_N_reg_17 : LNQD1BWP7T port map(EN => n_1651, D => n_1601, Q => new_N(17));
  new_N_reg_18 : LNQD1BWP7T port map(EN => n_1651, D => n_1600, Q => new_N(18));
  new_N_reg_19 : LNQD1BWP7T port map(EN => n_1651, D => n_1599, Q => new_N(19));
  new_N_reg_20 : LNQD1BWP7T port map(EN => n_1651, D => n_1598, Q => new_N(20));
  new_N_reg_21 : LNQD1BWP7T port map(EN => n_1651, D => n_1597, Q => new_N(21));
  new_N_reg_22 : LNQD1BWP7T port map(EN => n_1651, D => n_1596, Q => new_N(22));
  new_N_reg_23 : LNQD1BWP7T port map(EN => n_1651, D => n_1595, Q => new_N(23));
  new_N_reg_24 : LNQD1BWP7T port map(EN => n_1651, D => n_1594, Q => new_N(24));
  new_N_reg_25 : LNQD1BWP7T port map(EN => n_1651, D => n_1593, Q => new_N(25));
  new_N_reg_26 : LNQD1BWP7T port map(EN => n_1651, D => n_1592, Q => new_N(26));
  new_N_reg_27 : LNQD1BWP7T port map(EN => n_1651, D => n_1591, Q => new_N(27));
  new_N_reg_28 : LNQD1BWP7T port map(EN => n_1651, D => n_1590, Q => new_N(28));
  new_N_reg_29 : LNQD1BWP7T port map(EN => n_1651, D => n_1589, Q => new_N(29));
  new_N_reg_30 : LNQD1BWP7T port map(EN => n_1651, D => n_1588, Q => new_N(30));
  new_N_reg_31 : LNQD1BWP7T port map(EN => n_1651, D => n_1587, Q => new_N(31));
  new_corner_count_reg_1 : LHQD1BWP7T port map(E => n_1657, D => n_1648, Q => new_corner_count(1));
  new_corner_count_reg_2 : LHQD1BWP7T port map(E => n_1657, D => n_1647, Q => new_corner_count(2));
  new_corner_count_reg_3 : LHQD1BWP7T port map(E => n_1657, D => n_1646, Q => new_corner_count(3));
  new_corner_count_reg_4 : LHQD1BWP7T port map(E => n_1657, D => n_1645, Q => new_corner_count(4));
  new_corner_count_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1644, Q => new_corner_count(5));
  new_corner_count_reg_6 : LHQD1BWP7T port map(E => n_1657, D => n_1643, Q => new_corner_count(6));
  new_corner_count_reg_7 : LHQD1BWP7T port map(E => n_1657, D => n_1642, Q => new_corner_count(7));
  new_corner_count_reg_8 : LHQD1BWP7T port map(E => n_1657, D => n_1641, Q => new_corner_count(8));
  new_corner_count_reg_9 : LHQD1BWP7T port map(E => n_1657, D => n_1640, Q => new_corner_count(9));
  new_corner_count_reg_10 : LHQD1BWP7T port map(E => n_1657, D => n_1639, Q => new_corner_count(10));
  new_corner_count_reg_11 : LHQD1BWP7T port map(E => n_1657, D => n_1638, Q => new_corner_count(11));
  new_corner_count_reg_12 : LHQD1BWP7T port map(E => n_1657, D => n_1637, Q => new_corner_count(12));
  new_corner_count_reg_13 : LHQD1BWP7T port map(E => n_1657, D => n_1636, Q => new_corner_count(13));
  new_corner_count_reg_14 : LHQD1BWP7T port map(E => n_1657, D => n_1635, Q => new_corner_count(14));
  new_corner_count_reg_15 : LHQD1BWP7T port map(E => n_1657, D => n_1634, Q => new_corner_count(15));
  new_corner_count_reg_16 : LHQD1BWP7T port map(E => n_1657, D => n_1633, Q => new_corner_count(16));
  new_corner_count_reg_17 : LHQD1BWP7T port map(E => n_1657, D => n_1632, Q => new_corner_count(17));
  new_corner_count_reg_18 : LHQD1BWP7T port map(E => n_1657, D => n_1631, Q => new_corner_count(18));
  new_corner_count_reg_19 : LHQD1BWP7T port map(E => n_1657, D => n_1630, Q => new_corner_count(19));
  new_corner_count_reg_20 : LHQD1BWP7T port map(E => n_1657, D => n_1629, Q => new_corner_count(20));
  new_corner_count_reg_21 : LHQD1BWP7T port map(E => n_1657, D => n_1628, Q => new_corner_count(21));
  new_corner_count_reg_22 : LHQD1BWP7T port map(E => n_1657, D => n_1627, Q => new_corner_count(22));
  new_corner_count_reg_23 : LHQD1BWP7T port map(E => n_1657, D => n_1626, Q => new_corner_count(23));
  new_corner_count_reg_24 : LHQD1BWP7T port map(E => n_1657, D => n_1625, Q => new_corner_count(24));
  new_corner_count_reg_25 : LHQD1BWP7T port map(E => n_1657, D => n_1624, Q => new_corner_count(25));
  new_corner_count_reg_26 : LHQD1BWP7T port map(E => n_1657, D => n_1623, Q => new_corner_count(26));
  new_corner_count_reg_27 : LHQD1BWP7T port map(E => n_1657, D => n_1622, Q => new_corner_count(27));
  new_corner_count_reg_28 : LHQD1BWP7T port map(E => n_1657, D => n_1621, Q => new_corner_count(28));
  new_corner_count_reg_29 : LHQD1BWP7T port map(E => n_1657, D => n_1620, Q => new_corner_count(29));
  new_corner_count_reg_30 : LHQD1BWP7T port map(E => n_1657, D => n_1619, Q => new_corner_count(30));
  new_corner_count_reg_31 : LHQD1BWP7T port map(E => n_1657, D => n_1618, Q => new_corner_count(31));
  new_state_reg_0 : LHQD1BWP7T port map(E => n_1649, D => n_1040, Q => new_state(0));
  new_state_reg_1 : LHQD1BWP7T port map(E => n_1649, D => n_1041, Q => new_state(1));
  shift0_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output0(0), Q => shift0(0));
  shift0_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output0(1), Q => shift0(1));
  shift0_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output0(2), Q => shift0(2));
  shift0_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output0(3), Q => shift0(3));
  shift0_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output0(4), Q => shift0(4));
  shift0_reg_5 : LHQD1BWP7T port map(E => n_1657, D => snake_output0(5), Q => shift0(5));
  shift1_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output1(0), Q => shift1(0));
  shift1_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output1(1), Q => shift1(1));
  shift1_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output1(2), Q => shift1(2));
  shift1_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output1(3), Q => shift1(3));
  shift1_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output1(4), Q => shift1(4));
  shift1_reg_5 : LHQD1BWP7T port map(E => n_1657, D => snake_output1(5), Q => shift1(5));
  shift2_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output2(0), Q => shift2(0));
  shift2_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output2(1), Q => shift2(1));
  shift2_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output2(2), Q => shift2(2));
  shift2_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output2(3), Q => shift2(3));
  shift2_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output2(4), Q => shift2(4));
  shift2_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1179, Q => shift2(5));
  shift3_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output3(0), Q => shift3(0));
  shift3_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output3(1), Q => shift3(1));
  shift3_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output3(2), Q => shift3(2));
  shift3_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output3(3), Q => shift3(3));
  shift3_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output3(4), Q => shift3(4));
  shift3_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1173, Q => shift3(5));
  shift4_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output4(0), Q => shift4(0));
  shift4_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output4(1), Q => shift4(1));
  shift4_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output4(2), Q => shift4(2));
  shift4_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output4(3), Q => shift4(3));
  shift4_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output4(4), Q => shift4(4));
  shift4_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1167, Q => shift4(5));
  shift5_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output5(0), Q => shift5(0));
  shift5_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output5(1), Q => shift5(1));
  shift5_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output5(2), Q => shift5(2));
  shift5_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output5(3), Q => shift5(3));
  shift5_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output5(4), Q => shift5(4));
  shift5_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1161, Q => shift5(5));
  shift6_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output6(0), Q => shift6(0));
  shift6_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output6(1), Q => shift6(1));
  shift6_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output6(2), Q => shift6(2));
  shift6_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output6(3), Q => shift6(3));
  shift6_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output6(4), Q => shift6(4));
  shift6_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1155, Q => shift6(5));
  shift7_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output7(0), Q => shift7(0));
  shift7_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output7(1), Q => shift7(1));
  shift7_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output7(2), Q => shift7(2));
  shift7_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output7(3), Q => shift7(3));
  shift7_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output7(4), Q => shift7(4));
  shift7_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1149, Q => shift7(5));
  shift8_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output8(0), Q => shift8(0));
  shift8_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output8(1), Q => shift8(1));
  shift8_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output8(2), Q => shift8(2));
  shift8_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output8(3), Q => shift8(3));
  shift8_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output8(4), Q => shift8(4));
  shift8_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1143, Q => shift8(5));
  shift9_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output9(0), Q => shift9(0));
  shift9_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output9(1), Q => shift9(1));
  shift9_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output9(2), Q => shift9(2));
  shift9_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output9(3), Q => shift9(3));
  shift9_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output9(4), Q => shift9(4));
  shift9_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1137, Q => shift9(5));
  shift10_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output10(0), Q => shift10(0));
  shift10_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output10(1), Q => shift10(1));
  shift10_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output10(2), Q => shift10(2));
  shift10_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output10(3), Q => shift10(3));
  shift10_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output10(4), Q => shift10(4));
  shift10_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1131, Q => shift10(5));
  shift11_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output11(0), Q => shift11(0));
  shift11_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output11(1), Q => shift11(1));
  shift11_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output11(2), Q => shift11(2));
  shift11_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output11(3), Q => shift11(3));
  shift11_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output11(4), Q => shift11(4));
  shift11_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1125, Q => shift11(5));
  shift12_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output12(0), Q => shift12(0));
  shift12_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output12(1), Q => shift12(1));
  shift12_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output12(2), Q => shift12(2));
  shift12_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output12(3), Q => shift12(3));
  shift12_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output12(4), Q => shift12(4));
  shift12_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1119, Q => shift12(5));
  shift13_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output13(0), Q => shift13(0));
  shift13_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output13(1), Q => shift13(1));
  shift13_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output13(2), Q => shift13(2));
  shift13_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output13(3), Q => shift13(3));
  shift13_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output13(4), Q => shift13(4));
  shift13_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1113, Q => shift13(5));
  shift14_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output14(0), Q => shift14(0));
  shift14_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output14(1), Q => shift14(1));
  shift14_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output14(2), Q => shift14(2));
  shift14_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output14(3), Q => shift14(3));
  shift14_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output14(4), Q => shift14(4));
  shift14_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1107, Q => shift14(5));
  shift15_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output15(0), Q => shift15(0));
  shift15_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output15(1), Q => shift15(1));
  shift15_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output15(2), Q => shift15(2));
  shift15_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output15(3), Q => shift15(3));
  shift15_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output15(4), Q => shift15(4));
  shift15_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1101, Q => shift15(5));
  shift16_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output16(0), Q => shift16(0));
  shift16_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output16(1), Q => shift16(1));
  shift16_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output16(2), Q => shift16(2));
  shift16_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output16(3), Q => shift16(3));
  shift16_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output16(4), Q => shift16(4));
  shift16_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1095, Q => shift16(5));
  shift17_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output17(0), Q => shift17(0));
  shift17_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output17(1), Q => shift17(1));
  shift17_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output17(2), Q => shift17(2));
  shift17_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output17(3), Q => shift17(3));
  shift17_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output17(4), Q => shift17(4));
  shift17_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1089, Q => shift17(5));
  shift18_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output18(0), Q => shift18(0));
  shift18_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output18(1), Q => shift18(1));
  shift18_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output18(2), Q => shift18(2));
  shift18_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output18(3), Q => shift18(3));
  shift18_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output18(4), Q => shift18(4));
  shift18_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1083, Q => shift18(5));
  shift19_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output19(0), Q => shift19(0));
  shift19_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output19(1), Q => shift19(1));
  shift19_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output19(2), Q => shift19(2));
  shift19_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output19(3), Q => shift19(3));
  shift19_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output19(4), Q => shift19(4));
  shift19_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1077, Q => shift19(5));
  shift20_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output20(0), Q => shift20(0));
  shift20_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output20(1), Q => shift20(1));
  shift20_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output20(2), Q => shift20(2));
  shift20_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output20(3), Q => shift20(3));
  shift20_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output20(4), Q => shift20(4));
  shift20_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1071, Q => shift20(5));
  shift21_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output21(0), Q => shift21(0));
  shift21_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output21(1), Q => shift21(1));
  shift21_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output21(2), Q => shift21(2));
  shift21_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output21(3), Q => shift21(3));
  shift21_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output21(4), Q => shift21(4));
  shift21_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1065, Q => shift21(5));
  shift22_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output22(0), Q => shift22(0));
  shift22_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output22(1), Q => shift22(1));
  shift22_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output22(2), Q => shift22(2));
  shift22_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output22(3), Q => shift22(3));
  shift22_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output22(4), Q => shift22(4));
  shift22_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1059, Q => shift22(5));
  shift23_reg_0 : LHQD1BWP7T port map(E => n_1657, D => snake_output23(0), Q => shift23(0));
  shift23_reg_1 : LHQD1BWP7T port map(E => n_1657, D => snake_output23(1), Q => shift23(1));
  shift23_reg_2 : LHQD1BWP7T port map(E => n_1657, D => snake_output23(2), Q => shift23(2));
  shift23_reg_3 : LHQD1BWP7T port map(E => n_1657, D => snake_output23(3), Q => shift23(3));
  shift23_reg_4 : LHQD1BWP7T port map(E => n_1657, D => snake_output23(4), Q => shift23(4));
  shift23_reg_5 : LHQD1BWP7T port map(E => n_1657, D => n_1053, Q => shift23(5));
  snake_list_reg_1 : LHQD1BWP7T port map(E => n_1652, D => n_992, Q => n_1186);
  snake_list_reg_2 : LHQD1BWP7T port map(E => n_1652, D => n_991, Q => n_1187);
  snake_list_reg_3 : LHQD1BWP7T port map(E => n_1652, D => n_990, Q => n_1188);
  snake_list_reg_4 : LHQD1BWP7T port map(E => n_1652, D => n_989, Q => n_1189);
  snake_list_reg_5 : LHQD1BWP7T port map(E => n_1652, D => n_988, Q => n_1190);
  snake_list_reg_6 : LHQD1BWP7T port map(E => n_1652, D => n_952, Q => n_1191);
  snake_list_reg_7 : LHQD1BWP7T port map(E => n_1652, D => n_1018, Q => n_1192);
  snake_list_reg_8 : LHQD1BWP7T port map(E => n_1652, D => n_1030, Q => n_1193);
  snake_list_reg_9 : LHQD1BWP7T port map(E => n_1652, D => n_1017, Q => n_1194);
  snake_list_reg_10 : LHQD1BWP7T port map(E => n_1652, D => n_1023, Q => n_1195);
  snake_list_reg_11 : LHQD1BWP7T port map(E => n_1652, D => n_1029, Q => n_1196);
  snake_list_reg_12 : LHQD1BWP7T port map(E => n_1652, D => n_1028, Q => n_1197);
  snake_list_reg_13 : LHQD1BWP7T port map(E => n_1652, D => n_1026, Q => n_1198);
  snake_list_reg_14 : LHQD1BWP7T port map(E => n_1652, D => n_1016, Q => n_1199);
  snake_list_reg_15 : LHQD1BWP7T port map(E => n_1652, D => n_1031, Q => n_1200);
  snake_list_reg_16 : LHQD1BWP7T port map(E => n_1652, D => n_1025, Q => n_1201);
  state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => new_state(1), D => n_157, Q => state(1));
  state_reg_3 : DFKCNQD1BWP7T port map(CP => clk, CN => new_state(3), D => n_157, Q => state(3));
  state_reg_4 : DFKCNQD1BWP7T port map(CP => clk, CN => new_state(4), D => n_157, Q => state(4));
  g29160 : OR4D0BWP7T port map(A1 => n_1736, A2 => n_1748, A3 => n_236, A4 => n_1039, Z => n_1041);
  g29161 : NR4D0BWP7T port map(A1 => n_1039, A2 => n_236, A3 => n_676, A4 => n_1657, ZN => n_1040);
  g29162 : NR3D0BWP7T port map(A1 => n_1032, A2 => n_1038, A3 => n_1022, ZN => n_1039);
  g29164 : AO211D0BWP7T port map(A1 => n_1036, A2 => n_419, B => n_1035, C => n_1021, Z => n_1038);
  g29165 : OAI211D0BWP7T port map(A1 => n_221, A2 => n_472, B => n_1034, C => n_494, ZN => n_1037);
  g29166 : INR4D0BWP7T port map(A1 => n_1024, B1 => corner_count(11), B2 => corner_count(12), B3 => corner_count(4), ZN => n_1036);
  g29167 : OAI221D0BWP7T port map(A1 => n_1012, A2 => new_tail(2), B1 => new_tail(0), B2 => n_1013, C => n_1033, ZN => n_1035);
  g29168 : OA221D0BWP7T port map(A1 => n_473, A2 => n_213, B1 => n_440, B2 => n_471, C => n_1027, Z => n_1034);
  g29176 : AOI221D0BWP7T port map(A1 => n_1012, A2 => new_tail(2), B1 => n_1013, B2 => new_tail(0), C => n_1020, ZN => n_1033);
  g29177 : OAI211D0BWP7T port map(A1 => new_tail(4), A2 => n_1015, B => n_1571, C => n_1019, ZN => n_1032);
  g29178 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_984, B => n_1003, C => n_456, ZN => n_1031);
  g29181 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_995, B => n_1007, C => n_444, ZN => n_1030);
  g29182 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_987, B => n_1002, C => n_450, ZN => n_1029);
  g29183 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_976, B => n_1001, C => n_454, ZN => n_1028);
  g29185 : AN4D1BWP7T port map(A1 => n_1000, A2 => n_679, A3 => n_526, A4 => n_490, Z => n_1027);
  g29186 : OAI211D0BWP7T port map(A1 => n_203, A2 => n_995, B => n_1005, C => n_455, ZN => n_1026);
  g29187 : OAI211D0BWP7T port map(A1 => n_203, A2 => n_987, B => n_1004, C => n_459, ZN => n_1025);
  g29188 : INR4D0BWP7T port map(A1 => n_999, B1 => corner_count(8), B2 => corner_count(9), B3 => corner_count(10), ZN => n_1024);
  g29189 : OAI211D0BWP7T port map(A1 => n_203, A2 => n_984, B => n_1006, C => n_447, ZN => n_1023);
  g29190 : MOAI22D0BWP7T port map(A1 => n_1008, A2 => new_tail(5), B1 => n_1008, B2 => new_tail(5), ZN => n_1022);
  g29191 : MOAI22D0BWP7T port map(A1 => n_1014, A2 => new_tail(3), B1 => n_1014, B2 => new_tail(3), ZN => n_1021);
  g29192 : MOAI22D0BWP7T port map(A1 => n_1011, A2 => new_tail(1), B1 => n_1011, B2 => new_tail(1), ZN => n_1020);
  g29193 : ND2D0BWP7T port map(A1 => n_1015, A2 => new_tail(4), ZN => n_1019);
  g29194 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_994, B => n_998, C => n_443, ZN => n_1018);
  g29195 : OAI221D0BWP7T port map(A1 => n_985, A2 => n_203, B1 => n_155, B2 => n_208, C => n_1009, ZN => n_1017);
  g29196 : OAI221D0BWP7T port map(A1 => n_997, A2 => n_203, B1 => n_155, B2 => n_206, C => n_1010, ZN => n_1016);
  g29197 : OA21D0BWP7T port map(A1 => n_985, A2 => n_205, B => n_453, Z => n_1010);
  g29198 : OA21D0BWP7T port map(A1 => n_997, A2 => n_205, B => n_445, Z => n_1009);
  g29199 : AN4D1BWP7T port map(A1 => n_977, A2 => n_786, A3 => n_787, A4 => n_743, Z => n_1015);
  g29200 : AN4D1BWP7T port map(A1 => n_978, A2 => n_783, A3 => n_784, A4 => n_744, Z => n_1014);
  g29201 : AN4D1BWP7T port map(A1 => n_979, A2 => n_780, A3 => n_781, A4 => n_745, Z => n_1013);
  g29202 : AN4D1BWP7T port map(A1 => n_980, A2 => n_777, A3 => n_778, A4 => n_746, Z => n_1012);
  g29203 : AN4D1BWP7T port map(A1 => n_981, A2 => n_774, A3 => n_775, A4 => n_747, Z => n_1011);
  g29204 : AOI22D0BWP7T port map(A1 => n_996, A2 => n_202, B1 => n_1737, B2 => head(1), ZN => n_1007);
  g29205 : AOI22D0BWP7T port map(A1 => n_983, A2 => n_204, B1 => n_1737, B2 => head(3), ZN => n_1006);
  g29206 : AOI22D0BWP7T port map(A1 => n_996, A2 => n_204, B1 => n_1737, B2 => head(6), ZN => n_1005);
  g29207 : AOI22D0BWP7T port map(A1 => n_986, A2 => n_204, B1 => n_1737, B2 => head(9), ZN => n_1004);
  g29208 : AOI22D0BWP7T port map(A1 => n_983, A2 => n_202, B1 => n_1737, B2 => head(8), ZN => n_1003);
  g29209 : AOI22D0BWP7T port map(A1 => n_986, A2 => n_202, B1 => n_1737, B2 => head(4), ZN => n_1002);
  g29210 : MAOI22D0BWP7T port map(A1 => n_1737, A2 => head(5), B1 => n_994, B2 => n_203, ZN => n_1001);
  g29211 : AN4D1BWP7T port map(A1 => n_982, A2 => n_790, A3 => n_791, A4 => n_717, Z => n_1008);
  g29216 : AOI21D0BWP7T port map(A1 => n_1735, A2 => snake_output1(5), B => n_993, ZN => n_1000);
  g29217 : INR4D0BWP7T port map(A1 => n_969, B1 => corner_count(5), B2 => corner_count(6), B3 => corner_count(7), ZN => n_999);
  g29219 : MAOI22D0BWP7T port map(A1 => n_1737, A2 => head(0), B1 => n_976, B2 => n_203, ZN => n_998);
  g29220 : OAI21D0BWP7T port map(A1 => n_599, A2 => n_230, B => n_975, ZN => n_993);
  g29221 : ND4D0BWP7T port map(A1 => n_966, A2 => n_818, A3 => n_819, A4 => n_730, ZN => n_992);
  g29222 : ND4D0BWP7T port map(A1 => n_965, A2 => n_815, A3 => n_816, A4 => n_729, ZN => n_991);
  g29223 : ND4D0BWP7T port map(A1 => n_964, A2 => n_813, A3 => n_820, A4 => n_726, ZN => n_990);
  g29224 : ND4D0BWP7T port map(A1 => n_957, A2 => n_828, A3 => n_827, A4 => n_724, ZN => n_989);
  g29225 : ND4D0BWP7T port map(A1 => n_962, A2 => n_831, A3 => n_830, A4 => n_722, ZN => n_988);
  g29226 : AN4D1BWP7T port map(A1 => n_958, A2 => n_711, A3 => n_654, A4 => n_655, Z => n_997);
  g29227 : ND4D0BWP7T port map(A1 => n_959, A2 => n_713, A3 => n_586, A4 => n_658, ZN => n_996);
  g29228 : AN4D1BWP7T port map(A1 => n_960, A2 => n_715, A3 => n_665, A4 => n_666, Z => n_995);
  g29229 : AN4D1BWP7T port map(A1 => n_961, A2 => n_720, A3 => n_624, A4 => n_678, Z => n_994);
  g29230 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(5), B1 => n_605, B2 => snake_output21(5), C => n_972, ZN => n_982);
  g29231 : AOI221D0BWP7T port map(A1 => n_0, A2 => n_1091, B1 => n_605, B2 => n_1061, C => n_967, ZN => n_981);
  g29232 : AOI221D0BWP7T port map(A1 => n_0, A2 => n_1092, B1 => n_605, B2 => n_1062, C => n_968, ZN => n_980);
  g29233 : AOI221D0BWP7T port map(A1 => n_0, A2 => n_1090, B1 => n_605, B2 => n_1060, C => n_974, ZN => n_979);
  g29234 : AOI221D0BWP7T port map(A1 => n_0, A2 => n_1093, B1 => n_605, B2 => n_1063, C => n_970, ZN => n_978);
  g29235 : AOI221D0BWP7T port map(A1 => n_0, A2 => n_1094, B1 => n_605, B2 => n_1064, C => n_971, ZN => n_977);
  g29236 : AN4D1BWP7T port map(A1 => n_954, A2 => n_705, A3 => n_638, A4 => n_639, Z => n_987);
  g29237 : ND4D0BWP7T port map(A1 => n_953, A2 => n_704, A3 => n_576, A4 => n_634, ZN => n_986);
  g29238 : AN4D1BWP7T port map(A1 => n_963, A2 => n_710, A3 => n_582, A4 => n_649, Z => n_985);
  g29239 : AN4D1BWP7T port map(A1 => n_955, A2 => n_707, A3 => n_579, A4 => n_642, Z => n_984);
  g29240 : ND4D0BWP7T port map(A1 => n_956, A2 => n_708, A3 => n_645, A4 => n_646, ZN => n_983);
  g29242 : AOI31D0BWP7T port map(A1 => n_427, A2 => n_226, A3 => n_1113, B => n_973, ZN => n_975);
  g29243 : AN4D1BWP7T port map(A1 => n_951, A2 => n_719, A3 => n_589, A4 => n_668, Z => n_976);
  g29244 : ND4D0BWP7T port map(A1 => n_947, A2 => n_735, A3 => n_568, A4 => n_567, ZN => n_974);
  g29245 : IOA21D0BWP7T port map(A1 => n_940, A2 => n_1736, B => n_822, ZN => n_973);
  g29246 : ND4D0BWP7T port map(A1 => n_950, A2 => n_731, A3 => n_574, A4 => n_573, ZN => n_972);
  g29247 : ND4D0BWP7T port map(A1 => n_949, A2 => n_732, A3 => n_571, A4 => n_572, ZN => n_971);
  g29248 : ND4D0BWP7T port map(A1 => n_948, A2 => n_733, A3 => n_569, A4 => n_570, ZN => n_970);
  g29249 : INR4D0BWP7T port map(A1 => n_927, B1 => corner_count(19), B2 => corner_count(17), B3 => corner_count(18), ZN => n_969);
  g29250 : ND4D0BWP7T port map(A1 => n_946, A2 => n_736, A3 => n_591, A4 => n_578, ZN => n_968);
  g29251 : ND4D0BWP7T port map(A1 => n_945, A2 => n_737, A3 => n_593, A4 => n_592, ZN => n_967);
  g29252 : AOI221D0BWP7T port map(A1 => n_465, A2 => n_1096, B1 => n_560, B2 => n_1060, C => n_944, ZN => n_966);
  g29253 : AOI221D0BWP7T port map(A1 => n_465, A2 => n_1097, B1 => n_560, B2 => n_1061, C => n_943, ZN => n_965);
  g29254 : AOI221D0BWP7T port map(A1 => n_465, A2 => n_1098, B1 => n_560, B2 => n_1062, C => n_942, ZN => n_964);
  g29255 : AOI221D0BWP7T port map(A1 => n_562, A2 => n_1050, B1 => n_534, B2 => n_1080, C => n_938, ZN => n_963);
  g29256 : AOI221D0BWP7T port map(A1 => n_465, A2 => n_1100, B1 => n_560, B2 => n_1064, C => n_935, ZN => n_962);
  g29257 : AOI221D0BWP7T port map(A1 => n_515, A2 => n_1084, B1 => n_602, B2 => n_1054, C => n_934, ZN => n_961);
  g29258 : AOI221D0BWP7T port map(A1 => n_515, A2 => n_1085, B1 => n_602, B2 => n_1055, C => n_933, ZN => n_960);
  g29259 : AOI221D0BWP7T port map(A1 => n_562, A2 => n_1049, B1 => n_534, B2 => n_1079, C => n_939, ZN => n_959);
  g29260 : AOI221D0BWP7T port map(A1 => n_515, A2 => n_1086, B1 => n_602, B2 => n_1056, C => n_932, ZN => n_958);
  g29261 : AOI221D0BWP7T port map(A1 => n_465, A2 => n_1099, B1 => n_560, B2 => n_1063, C => n_941, ZN => n_957);
  g29262 : AOI221D0BWP7T port map(A1 => n_515, A2 => n_1087, B1 => n_602, B2 => n_1057, C => n_931, ZN => n_956);
  g29263 : AOI221D0BWP7T port map(A1 => n_562, A2 => n_1051, B1 => n_534, B2 => n_1081, C => n_937, ZN => n_955);
  g29264 : AOI221D0BWP7T port map(A1 => n_515, A2 => n_1088, B1 => n_602, B2 => n_1058, C => n_930, ZN => n_954);
  g29265 : AOI221D0BWP7T port map(A1 => n_562, A2 => n_1052, B1 => n_534, B2 => n_1082, C => n_936, ZN => n_953);
  g29266 : AO22D0BWP7T port map(A1 => n_940, A2 => n_192, B1 => snake_output0(5), B2 => n_1737, Z => n_952);
  g29267 : AOI221D0BWP7T port map(A1 => n_562, A2 => n_1048, B1 => n_534, B2 => n_1078, C => n_922, ZN => n_951);
  g29268 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(5), B1 => n_518, B2 => snake_output15(5), C => n_928, ZN => n_950);
  g29269 : AOI221D0BWP7T port map(A1 => n_517, A2 => n_1106, B1 => n_518, B2 => n_1100, C => n_929, ZN => n_949);
  g29270 : AOI221D0BWP7T port map(A1 => n_517, A2 => n_1105, B1 => n_518, B2 => n_1099, C => n_926, ZN => n_948);
  g29271 : AOI221D0BWP7T port map(A1 => n_517, A2 => n_1102, B1 => n_518, B2 => n_1096, C => n_923, ZN => n_947);
  g29272 : AOI221D0BWP7T port map(A1 => n_517, A2 => n_1104, B1 => n_518, B2 => n_1098, C => n_924, ZN => n_946);
  g29273 : AOI221D0BWP7T port map(A1 => n_517, A2 => n_1103, B1 => n_518, B2 => n_1097, C => n_925, ZN => n_945);
  g29274 : ND4D0BWP7T port map(A1 => n_906, A2 => n_861, A3 => n_853, A4 => n_680, ZN => n_944);
  g29275 : ND4D0BWP7T port map(A1 => n_910, A2 => n_826, A3 => n_728, A4 => n_814, ZN => n_943);
  g29276 : ND4D0BWP7T port map(A1 => n_909, A2 => n_825, A3 => n_852, A4 => n_821, ZN => n_942);
  g29277 : ND4D0BWP7T port map(A1 => n_908, A2 => n_824, A3 => n_851, A4 => n_829, ZN => n_941);
  g29278 : ND4D0BWP7T port map(A1 => n_916, A2 => n_712, A3 => n_657, A4 => n_628, ZN => n_939);
  g29279 : ND4D0BWP7T port map(A1 => n_915, A2 => n_709, A3 => n_648, A4 => n_627, ZN => n_938);
  g29280 : ND4D0BWP7T port map(A1 => n_914, A2 => n_706, A3 => n_641, A4 => n_626, ZN => n_937);
  g29281 : ND4D0BWP7T port map(A1 => n_913, A2 => n_703, A3 => n_633, A4 => n_625, ZN => n_936);
  g29282 : ND4D0BWP7T port map(A1 => n_907, A2 => n_823, A3 => n_850, A4 => n_832, ZN => n_935);
  g29283 : ND4D0BWP7T port map(A1 => n_921, A2 => n_671, A3 => n_833, A4 => n_834, ZN => n_934);
  g29284 : ND4D0BWP7T port map(A1 => n_920, A2 => n_663, A3 => n_838, A4 => n_839, ZN => n_933);
  g29285 : ND4D0BWP7T port map(A1 => n_919, A2 => n_653, A3 => n_806, A4 => n_805, ZN => n_932);
  g29286 : ND4D0BWP7T port map(A1 => n_918, A2 => n_644, A3 => n_801, A4 => n_800, ZN => n_931);
  g29287 : ND4D0BWP7T port map(A1 => n_917, A2 => n_637, A3 => n_796, A4 => n_795, ZN => n_930);
  g29288 : ND4D0BWP7T port map(A1 => n_912, A2 => n_718, A3 => n_716, A4 => n_672, ZN => n_940);
  g29289 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(4), B => n_911, Z => n_929);
  g29290 : AO21D0BWP7T port map(A1 => n_604, A2 => n_1047, B => n_901, Z => n_928);
  g29291 : INR4D0BWP7T port map(A1 => n_885, B1 => corner_count(22), B2 => corner_count(21), B3 => corner_count(20), ZN => n_927);
  g29292 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(3), B => n_905, Z => n_926);
  g29293 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(1), B => n_902, Z => n_925);
  g29294 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(2), B => n_903, Z => n_924);
  g29295 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(0), B => n_904, Z => n_923);
  g29296 : ND4D0BWP7T port map(A1 => n_898, A2 => n_837, A3 => n_836, A4 => n_588, ZN => n_922);
  g29297 : AOI221D0BWP7T port map(A1 => n_498, A2 => n_1168, B1 => n_510, B2 => n_1174, C => n_899, ZN => n_921);
  g29298 : AOI221D0BWP7T port map(A1 => n_498, A2 => n_1169, B1 => n_510, B2 => n_1175, C => n_900, ZN => n_920);
  g29299 : AOI221D0BWP7T port map(A1 => n_498, A2 => n_1170, B1 => n_510, B2 => n_1176, C => n_896, ZN => n_919);
  g29300 : AOI221D0BWP7T port map(A1 => n_498, A2 => n_1171, B1 => n_510, B2 => n_1177, C => n_894, ZN => n_918);
  g29301 : AOI221D0BWP7T port map(A1 => n_498, A2 => n_1172, B1 => n_510, B2 => n_1178, C => n_892, ZN => n_917);
  g29302 : AOI221D0BWP7T port map(A1 => n_475, A2 => snake_output14(1), B1 => n_418, B2 => n_1109, C => n_897, ZN => n_916);
  g29303 : AOI221D0BWP7T port map(A1 => n_514, A2 => n_1122, B1 => n_475, B2 => n_1104, C => n_893, ZN => n_915);
  g29304 : AOI221D0BWP7T port map(A1 => n_514, A2 => n_1123, B1 => n_475, B2 => n_1105, C => n_895, ZN => n_914);
  g29305 : AOI221D0BWP7T port map(A1 => n_514, A2 => n_1124, B1 => n_475, B2 => n_1106, C => n_891, ZN => n_913);
  g29306 : NR3D0BWP7T port map(A1 => n_869, A2 => n_871, A3 => n_810, ZN => n_912);
  g29307 : ND4D0BWP7T port map(A1 => n_877, A2 => n_848, A3 => n_785, A4 => n_772, ZN => n_911);
  g29308 : AOI221D0BWP7T port map(A1 => n_752, A2 => n_1139, B1 => n_480, B2 => n_1055, C => n_883, ZN => n_910);
  g29309 : AOI221D0BWP7T port map(A1 => n_618, A2 => n_1128, B1 => n_480, B2 => n_1056, C => n_882, ZN => n_909);
  g29310 : AOI221D0BWP7T port map(A1 => n_618, A2 => n_1129, B1 => n_480, B2 => n_1057, C => n_881, ZN => n_908);
  g29311 : AOI221D0BWP7T port map(A1 => n_618, A2 => n_1130, B1 => n_480, B2 => n_1058, C => n_880, ZN => n_907);
  g29312 : AOI221D0BWP7T port map(A1 => n_618, A2 => n_1126, B1 => n_480, B2 => n_1054, C => n_884, ZN => n_906);
  g29313 : ND4D0BWP7T port map(A1 => n_876, A2 => n_847, A3 => n_782, A4 => n_771, ZN => n_905);
  g29314 : ND4D0BWP7T port map(A1 => n_875, A2 => n_846, A3 => n_779, A4 => n_770, ZN => n_904);
  g29315 : ND4D0BWP7T port map(A1 => n_874, A2 => n_845, A3 => n_776, A4 => n_769, ZN => n_903);
  g29316 : ND4D0BWP7T port map(A1 => n_873, A2 => n_844, A3 => n_773, A4 => n_768, ZN => n_902);
  g29317 : ND4D0BWP7T port map(A1 => n_878, A2 => n_849, A3 => n_788, A4 => n_789, ZN => n_901);
  g29318 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(1), B => n_870, Z => n_900);
  g29319 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(0), B => n_872, Z => n_899);
  g29320 : AOI221D0BWP7T port map(A1 => n_510, A2 => n_1180, B1 => n_532, B2 => n_1156, C => n_879, ZN => n_898);
  g29321 : AO21D0BWP7T port map(A1 => n_621, A2 => n_1043, B => n_868, Z => n_897);
  g29322 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(2), B => n_867, Z => n_896);
  g29323 : AO21D0BWP7T port map(A1 => n_621, A2 => snake_output24(3), B => n_864, Z => n_895);
  g29324 : AO21D0BWP7T port map(A1 => n_611, A2 => n_1045, B => n_865, Z => n_894);
  g29325 : AO21D0BWP7T port map(A1 => n_621, A2 => n_1044, B => n_866, Z => n_893);
  g29326 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(4), B => n_863, Z => n_892);
  g29327 : AO21D0BWP7T port map(A1 => n_621, A2 => n_1046, B => n_862, Z => n_891);
  g29355 : INR4D0BWP7T port map(A1 => n_734, B1 => corner_count(25), B2 => corner_count(24), B3 => corner_count(23), ZN => n_885);
  g29356 : ND3D0BWP7T port map(A1 => n_843, A2 => n_738, A3 => n_681, ZN => n_884);
  g29357 : ND3D0BWP7T port map(A1 => n_857, A2 => n_739, A3 => n_682, ZN => n_883);
  g29358 : ND3D0BWP7T port map(A1 => n_856, A2 => n_740, A3 => n_683, ZN => n_882);
  g29359 : ND3D0BWP7T port map(A1 => n_855, A2 => n_741, A3 => n_677, ZN => n_881);
  g29360 : ND3D0BWP7T port map(A1 => n_854, A2 => n_742, A3 => n_675, ZN => n_880);
  g29361 : AO21D0BWP7T port map(A1 => n_621, A2 => n_1042, B => n_858, Z => n_879);
  g29362 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(5), B1 => n_841, B2 => snake_output7(5), ZN => n_878);
  g29363 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(4), B1 => n_841, B2 => n_1148, ZN => n_877);
  g29364 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(3), B1 => n_841, B2 => n_1147, ZN => n_876);
  g29365 : AOI22D0BWP7T port map(A1 => n_842, A2 => n_1150, B1 => n_841, B2 => n_1144, ZN => n_875);
  g29366 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(2), B1 => n_841, B2 => n_1146, ZN => n_874);
  g29367 : AOI22D0BWP7T port map(A1 => n_842, A2 => n_1151, B1 => n_841, B2 => n_1145, ZN => n_873);
  g29368 : ND4D0BWP7T port map(A1 => n_835, A2 => n_670, A3 => n_669, A4 => n_590, ZN => n_872);
  g29369 : ND4D0BWP7T port map(A1 => n_808, A2 => n_662, A3 => n_660, A4 => n_714, ZN => n_871);
  g29370 : ND4D0BWP7T port map(A1 => n_840, A2 => n_661, A3 => n_659, A4 => n_587, ZN => n_870);
  g29371 : ND4D0BWP7T port map(A1 => n_652, A2 => n_584, A3 => n_807, A4 => n_630, ZN => n_869);
  g29372 : ND4D0BWP7T port map(A1 => n_809, A2 => n_767, A3 => n_585, A4 => n_656, ZN => n_868);
  g29373 : ND4D0BWP7T port map(A1 => n_804, A2 => n_651, A3 => n_650, A4 => n_583, ZN => n_867);
  g29374 : ND4D0BWP7T port map(A1 => n_803, A2 => n_802, A3 => n_581, A4 => n_647, ZN => n_866);
  g29375 : ND4D0BWP7T port map(A1 => n_799, A2 => n_632, A3 => n_643, A4 => n_580, ZN => n_865);
  g29376 : ND4D0BWP7T port map(A1 => n_797, A2 => n_594, A3 => n_798, A4 => n_640, ZN => n_864);
  g29377 : ND4D0BWP7T port map(A1 => n_794, A2 => n_636, A3 => n_635, A4 => n_577, ZN => n_863);
  g29378 : ND4D0BWP7T port map(A1 => n_792, A2 => n_793, A3 => n_575, A4 => n_631, ZN => n_862);
  g29382 : AOI221D0BWP7T port map(A1 => n_538, A2 => n_1090, B1 => n_558, B2 => n_1108, C => n_817, ZN => n_861);
  g29395 : OAI21D0BWP7T port map(A1 => n_1, A2 => n_1701, B => n_195, ZN => n_890);
  g29396 : AOI21D0BWP7T port map(A1 => n_754, A2 => n_222, B => n_194, ZN => n_886);
  g29397 : AOI21D0BWP7T port map(A1 => n_754, A2 => n_212, B => n_194, ZN => n_887);
  g29398 : OAI21D0BWP7T port map(A1 => n_753, A2 => n_217, B => n_195, ZN => n_889);
  g29399 : ND4D0BWP7T port map(A1 => n_748, A2 => n_667, A3 => n_629, A4 => n_527, ZN => n_858);
  g29400 : AOI222D0BWP7T port map(A1 => n_614, A2 => n_1181, B1 => n_616, B2 => n_1103, C1 => n_751, C2 => n_1157, ZN => n_857);
  g29401 : AOI222D0BWP7T port map(A1 => n_614, A2 => n_1182, B1 => n_616, B2 => n_1104, C1 => n_751, C2 => n_1158, ZN => n_856);
  g29402 : AOI222D0BWP7T port map(A1 => n_614, A2 => n_1183, B1 => n_616, B2 => n_1105, C1 => n_751, C2 => n_1159, ZN => n_855);
  g29403 : AOI222D0BWP7T port map(A1 => n_614, A2 => n_1184, B1 => n_616, B2 => n_1106, C1 => n_751, C2 => n_1160, ZN => n_854);
  g29404 : AOI22D0BWP7T port map(A1 => n_752, A2 => n_1138, B1 => n_615, B2 => n_1144, ZN => n_853);
  g29405 : AOI22D0BWP7T port map(A1 => n_752, A2 => n_1140, B1 => n_557, B2 => snake_output11(2), ZN => n_852);
  g29406 : AOI22D0BWP7T port map(A1 => n_752, A2 => n_1141, B1 => n_557, B2 => snake_output11(3), ZN => n_851);
  g29407 : AOI22D0BWP7T port map(A1 => n_752, A2 => n_1142, B1 => n_557, B2 => snake_output11(4), ZN => n_850);
  g29408 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(5), B1 => n_749, B2 => snake_output3(5), ZN => n_849);
  g29409 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(4), B1 => n_749, B2 => snake_output3(4), ZN => n_848);
  g29410 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(3), B1 => n_749, B2 => snake_output3(3), ZN => n_847);
  g29411 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(0), B1 => n_749, B2 => snake_output3(0), ZN => n_846);
  g29412 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(2), B1 => n_749, B2 => snake_output3(2), ZN => n_845);
  g29413 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(1), B1 => n_749, B2 => snake_output3(1), ZN => n_844);
  g29414 : AOI222D0BWP7T port map(A1 => n_614, A2 => n_1180, B1 => n_616, B2 => n_1102, C1 => n_751, C2 => n_1156, ZN => n_843);
  g29415 : OAI21D0BWP7T port map(A1 => n_753, A2 => n_220, B => n_195, ZN => n_888);
  g29416 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output8(1), B1 => n_554, B2 => n_1133, ZN => n_840);
  g29417 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1163, B1 => n_500, B2 => n_1157, ZN => n_839);
  g29418 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(1), B1 => n_532, B2 => snake_output6(1), ZN => n_838);
  g29419 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output7(0), B1 => n_685, B2 => n_1150, ZN => n_837);
  g29420 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1168, B1 => n_498, B2 => n_1174, ZN => n_836);
  g29421 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1138, B1 => n_554, B2 => snake_output9(0), ZN => n_835);
  g29422 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1162, B1 => n_500, B2 => n_1156, ZN => n_834);
  g29423 : AOI22D0BWP7T port map(A1 => n_685, A2 => n_1144, B1 => n_532, B2 => snake_output6(0), ZN => n_833);
  g29424 : AOI22D0BWP7T port map(A1 => n_698, A2 => n_1136, B1 => n_613, B2 => n_1118, ZN => n_832);
  g29425 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(4), B1 => n_697, B2 => snake_output23(4), ZN => n_831);
  g29426 : AOI22D0BWP7T port map(A1 => n_695, A2 => n_1076, B1 => n_696, B2 => n_1046, ZN => n_830);
  g29427 : AOI22D0BWP7T port map(A1 => n_698, A2 => n_1135, B1 => n_613, B2 => n_1117, ZN => n_829);
  g29428 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(3), B1 => n_697, B2 => snake_output23(3), ZN => n_828);
  g29429 : AOI22D0BWP7T port map(A1 => n_695, A2 => n_1075, B1 => n_696, B2 => n_1045, ZN => n_827);
  g29430 : AOI221D0BWP7T port map(A1 => n_561, A2 => n_1151, B1 => n_558, B2 => n_1109, C => n_727, ZN => n_826);
  g29431 : AOI221D0BWP7T port map(A1 => n_561, A2 => n_1152, B1 => n_558, B2 => n_1110, C => n_725, ZN => n_825);
  g29432 : AOI221D0BWP7T port map(A1 => n_561, A2 => n_1153, B1 => n_558, B2 => n_1111, C => n_723, ZN => n_824);
  g29433 : AOI221D0BWP7T port map(A1 => n_561, A2 => n_1154, B1 => n_558, B2 => n_1112, C => n_721, ZN => n_823);
  g29434 : OAI31D0BWP7T port map(A1 => n_600, A2 => n_1732, A3 => n_1737, B => snake_output0(5), ZN => n_822);
  g29435 : AOI22D0BWP7T port map(A1 => n_698, A2 => n_1134, B1 => n_613, B2 => n_1116, ZN => n_821);
  g29436 : AOI22D0BWP7T port map(A1 => n_695, A2 => n_1074, B1 => n_696, B2 => n_1044, ZN => n_820);
  g29437 : AOI22D0BWP7T port map(A1 => n_695, A2 => n_1072, B1 => n_696, B2 => n_1042, ZN => n_819);
  g29438 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(0), B1 => n_697, B2 => snake_output23(0), ZN => n_818);
  g29439 : AO22D0BWP7T port map(A1 => n_698, A2 => n_1132, B1 => n_1114, B2 => n_613, Z => n_817);
  g29440 : AOI22D0BWP7T port map(A1 => n_695, A2 => n_1073, B1 => n_696, B2 => n_1043, ZN => n_816);
  g29441 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(1), B1 => n_697, B2 => snake_output23(1), ZN => n_815);
  g29442 : AOI22D0BWP7T port map(A1 => n_698, A2 => n_1133, B1 => n_618, B2 => n_1127, ZN => n_814);
  g29443 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(2), B1 => n_697, B2 => snake_output23(2), ZN => n_813);
  g29446 : NR2D0BWP7T port map(A1 => n_755, A2 => corner_count(0), ZN => n_842);
  g29447 : NR2D0BWP7T port map(A1 => n_755, A2 => n_146, ZN => n_841);
  g29457 : AOI21D0BWP7T port map(A1 => n_700, A2 => n_1700, B => n_194, ZN => n_860);
  g29459 : OAI21D0BWP7T port map(A1 => n_701, A2 => n_1700, B => n_195, ZN => n_859);
  g29460 : MOAI22D0BWP7T port map(A1 => n_664, A2 => n_477, B1 => n_515, B2 => snake_output18(5), ZN => n_810);
  g29461 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1145, B1 => n_685, B2 => n_1151, ZN => n_809);
  g29462 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output8(5), B1 => n_554, B2 => snake_output10(5), ZN => n_808);
  g29463 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output5(5), B1 => n_496, B2 => snake_output2(5), ZN => n_807);
  g29464 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(2), B1 => n_532, B2 => n_1152, ZN => n_806);
  g29465 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1164, B1 => n_500, B2 => n_1158, ZN => n_805);
  g29466 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1140, B1 => n_554, B2 => n_1134, ZN => n_804);
  g29467 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1146, B1 => n_685, B2 => n_1152, ZN => n_803);
  g29468 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1170, B1 => n_498, B2 => n_1176, ZN => n_802);
  g29469 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(3), B1 => n_532, B2 => n_1153, ZN => n_801);
  g29470 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1165, B1 => n_500, B2 => n_1159, ZN => n_800);
  g29471 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1141, B1 => n_554, B2 => n_1135, ZN => n_799);
  g29472 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1171, B1 => n_496, B2 => snake_output0(3), ZN => n_798);
  g29473 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1147, B1 => n_685, B2 => n_1153, ZN => n_797);
  g29474 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(4), B1 => n_532, B2 => n_1154, ZN => n_796);
  g29475 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1166, B1 => n_500, B2 => n_1160, ZN => n_795);
  g29476 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1142, B1 => n_554, B2 => n_1136, ZN => n_794);
  g29477 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1172, B1 => n_498, B2 => n_1178, ZN => n_793);
  g29478 : AOI22D0BWP7T port map(A1 => n_688, A2 => n_1148, B1 => n_685, B2 => n_1154, ZN => n_792);
  g29479 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(5), B1 => n_606, B2 => snake_output18(5), ZN => n_791);
  g29480 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(5), B1 => n_608, B2 => snake_output17(5), ZN => n_790);
  g29481 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(5), B1 => n_693, B2 => snake_output5(5), ZN => n_789);
  g29482 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(5), B1 => n_689, B2 => n_1185, ZN => n_788);
  g29483 : AOI22D0BWP7T port map(A1 => n_692, A2 => n_1058, B1 => n_606, B2 => snake_output18(4), ZN => n_787);
  g29484 : AOI22D0BWP7T port map(A1 => n_691, A2 => n_1052, B1 => n_608, B2 => n_1088, ZN => n_786);
  g29485 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(4), B1 => n_689, B2 => n_1184, ZN => n_785);
  g29486 : AOI22D0BWP7T port map(A1 => n_692, A2 => n_1057, B1 => n_606, B2 => snake_output18(3), ZN => n_784);
  g29487 : AOI22D0BWP7T port map(A1 => n_691, A2 => n_1051, B1 => n_608, B2 => n_1087, ZN => n_783);
  g29488 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(3), B1 => n_689, B2 => n_1183, ZN => n_782);
  g29489 : AOI22D0BWP7T port map(A1 => n_692, A2 => n_1054, B1 => n_606, B2 => snake_output18(0), ZN => n_781);
  g29490 : AOI22D0BWP7T port map(A1 => n_691, A2 => n_1048, B1 => n_608, B2 => n_1084, ZN => n_780);
  g29491 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(0), B1 => n_689, B2 => n_1180, ZN => n_779);
  g29492 : AOI22D0BWP7T port map(A1 => n_692, A2 => n_1056, B1 => n_606, B2 => snake_output18(2), ZN => n_778);
  g29493 : AOI22D0BWP7T port map(A1 => n_691, A2 => n_1050, B1 => n_608, B2 => n_1086, ZN => n_777);
  g29494 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(2), B1 => n_689, B2 => n_1182, ZN => n_776);
  g29495 : AOI22D0BWP7T port map(A1 => n_692, A2 => n_1055, B1 => n_606, B2 => snake_output18(1), ZN => n_775);
  g29496 : AOI22D0BWP7T port map(A1 => n_691, A2 => n_1049, B1 => n_608, B2 => n_1085, ZN => n_774);
  g29497 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(1), B1 => n_689, B2 => n_1181, ZN => n_773);
  g29498 : AOI22D0BWP7T port map(A1 => n_690, A2 => n_1166, B1 => n_693, B2 => n_1160, ZN => n_772);
  g29499 : AOI22D0BWP7T port map(A1 => n_690, A2 => n_1165, B1 => n_693, B2 => n_1159, ZN => n_771);
  g29500 : AOI22D0BWP7T port map(A1 => n_690, A2 => n_1162, B1 => n_693, B2 => snake_output5(0), ZN => n_770);
  g29501 : AOI22D0BWP7T port map(A1 => n_690, A2 => n_1164, B1 => n_693, B2 => n_1158, ZN => n_769);
  g29502 : AOI22D0BWP7T port map(A1 => n_690, A2 => n_1163, B1 => n_693, B2 => n_1157, ZN => n_768);
  g29503 : AOI22D0BWP7T port map(A1 => n_687, A2 => n_1169, B1 => n_498, B2 => n_1175, ZN => n_767);
  g29567 : CKND1BWP7T port map(I => n_754, ZN => n_753);
  g29568 : AOI22D0BWP7T port map(A1 => n_617, A2 => snake_output8(0), B1 => n_512, B2 => n_1132, ZN => n_748);
  g29569 : AOI22D0BWP7T port map(A1 => n_607, A2 => n_1073, B1 => n_609, B2 => n_1067, ZN => n_747);
  g29570 : AOI22D0BWP7T port map(A1 => n_607, A2 => n_1074, B1 => n_609, B2 => n_1068, ZN => n_746);
  g29571 : AOI22D0BWP7T port map(A1 => n_607, A2 => n_1072, B1 => n_609, B2 => n_1066, ZN => n_745);
  g29572 : AOI22D0BWP7T port map(A1 => n_607, A2 => n_1075, B1 => n_609, B2 => n_1069, ZN => n_744);
  g29573 : AOI22D0BWP7T port map(A1 => n_607, A2 => n_1076, B1 => n_609, B2 => n_1070, ZN => n_743);
  g29574 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(4), B1 => n_537, B2 => n_1178, ZN => n_742);
  g29575 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(3), B1 => n_537, B2 => n_1177, ZN => n_741);
  g29576 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(2), B1 => n_537, B2 => n_1176, ZN => n_740);
  g29577 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(1), B1 => n_537, B2 => n_1175, ZN => n_739);
  g29578 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(0), B1 => n_537, B2 => n_1174, ZN => n_738);
  g29579 : AOI22D0BWP7T port map(A1 => n_603, A2 => n_1139, B1 => n_516, B2 => snake_output9(1), ZN => n_737);
  g29580 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(2), B1 => n_516, B2 => snake_output9(2), ZN => n_736);
  g29581 : AOI22D0BWP7T port map(A1 => n_603, A2 => n_1138, B1 => n_516, B2 => n_1132, ZN => n_735);
  g29582 : INR4D0BWP7T port map(A1 => n_528, B1 => corner_count(28), B2 => corner_count(27), B3 => corner_count(26), ZN => n_734);
  g29583 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(3), B1 => n_516, B2 => snake_output9(3), ZN => n_733);
  g29585 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(4), B1 => n_516, B2 => snake_output9(4), ZN => n_732);
  g29586 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(5), B1 => n_516, B2 => snake_output9(5), ZN => n_731);
  g29587 : AOI22D0BWP7T port map(A1 => n_612, A2 => n_1066, B1 => n_556, B2 => n_1078, ZN => n_730);
  g29588 : AOI22D0BWP7T port map(A1 => n_612, A2 => n_1067, B1 => n_556, B2 => n_1079, ZN => n_729);
  g29589 : AOI22D0BWP7T port map(A1 => n_557, A2 => n_1121, B1 => n_613, B2 => n_1115, ZN => n_728);
  g29590 : AO22D0BWP7T port map(A1 => n_538, A2 => n_1091, B1 => n_1145, B2 => n_615, Z => n_727);
  g29591 : AOI22D0BWP7T port map(A1 => n_612, A2 => n_1068, B1 => n_556, B2 => n_1080, ZN => n_726);
  g29592 : AO22D0BWP7T port map(A1 => n_538, A2 => n_1092, B1 => n_1146, B2 => n_615, Z => n_725);
  g29593 : AOI22D0BWP7T port map(A1 => n_612, A2 => n_1069, B1 => n_556, B2 => n_1081, ZN => n_724);
  g29594 : AO22D0BWP7T port map(A1 => n_538, A2 => n_1093, B1 => n_1147, B2 => n_615, Z => n_723);
  g29595 : AOI22D0BWP7T port map(A1 => n_612, A2 => n_1070, B1 => n_556, B2 => n_1082, ZN => n_722);
  g29596 : AO22D0BWP7T port map(A1 => n_538, A2 => n_1094, B1 => n_1148, B2 => n_615, Z => n_721);
  g29597 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1078, B1 => n_502, B2 => snake_output20(0), ZN => n_720);
  g29598 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1084, B1 => n_602, B2 => n_1060, ZN => n_719);
  g29599 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output19(5), B1 => n_534, B2 => snake_output20(5), ZN => n_718);
  g29600 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(5), B1 => n_609, B2 => snake_output20(5), ZN => n_717);
  g29601 : AOI22D0BWP7T port map(A1 => n_602, A2 => n_1053, B1 => n_502, B2 => n_1065, ZN => n_716);
  g29602 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1079, B1 => n_502, B2 => snake_output20(1), ZN => n_715);
  g29603 : AOI22D0BWP7T port map(A1 => n_622, A2 => n_1137, B1 => n_512, B2 => snake_output11(5), ZN => n_714);
  g29604 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1085, B1 => n_602, B2 => n_1061, ZN => n_713);
  g29605 : AOI22D0BWP7T port map(A1 => n_617, A2 => n_1139, B1 => n_512, B2 => n_1133, ZN => n_712);
  g29606 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1080, B1 => n_502, B2 => snake_output20(2), ZN => n_711);
  g29607 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1086, B1 => n_602, B2 => n_1062, ZN => n_710);
  g29608 : AOI22D0BWP7T port map(A1 => n_617, A2 => n_1140, B1 => n_512, B2 => n_1134, ZN => n_709);
  g29609 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1081, B1 => n_502, B2 => snake_output20(3), ZN => n_708);
  g29610 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1087, B1 => n_602, B2 => n_1063, ZN => n_707);
  g29611 : AOI22D0BWP7T port map(A1 => n_617, A2 => n_1141, B1 => n_512, B2 => n_1135, ZN => n_706);
  g29612 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1082, B1 => n_502, B2 => snake_output20(4), ZN => n_705);
  g29613 : AOI22D0BWP7T port map(A1 => n_596, A2 => n_1088, B1 => n_602, B2 => n_1064, ZN => n_704);
  g29614 : AOI22D0BWP7T port map(A1 => n_617, A2 => n_1142, B1 => n_512, B2 => n_1136, ZN => n_703);
  g29615 : ND2D0BWP7T port map(A1 => n_699, A2 => n_1740, ZN => n_755);
  g29616 : NR3D0BWP7T port map(A1 => n_610, A2 => n_1699, A3 => n_156, ZN => n_754);
  g29619 : NR2D0BWP7T port map(A1 => n_193, A2 => n_684, ZN => n_752);
  g29620 : NR2D0BWP7T port map(A1 => n_193, A2 => n_686, ZN => n_751);
  g29621 : OAI21D0BWP7T port map(A1 => n_610, A2 => n_434, B => n_195, ZN => n_811);
  g29622 : AN2D1BWP7T port map(A1 => n_699, A2 => n_231, Z => n_750);
  g29626 : AN2D1BWP7T port map(A1 => n_699, A2 => n_227, Z => n_749);
  g29631 : OAI21D0BWP7T port map(A1 => n_610, A2 => n_1581, B => n_195, ZN => n_812);
  g29632 : CKND1BWP7T port map(I => n_700, ZN => n_701);
  g29633 : INVD0BWP7T port map(I => n_687, ZN => n_686);
  g29634 : CKND1BWP7T port map(I => n_685, ZN => n_684);
  g29635 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(2), B1 => n_539, B2 => n_1170, ZN => n_683);
  g29636 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(1), B1 => n_539, B2 => n_1169, ZN => n_682);
  g29637 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(0), B1 => n_539, B2 => n_1168, ZN => n_681);
  g29638 : AOI22D0BWP7T port map(A1 => n_561, A2 => n_1150, B1 => n_557, B2 => n_1120, ZN => n_680);
  g29639 : AOI31D0BWP7T port map(A1 => n_1734, A2 => n_532, A3 => n_1143, B => n_547, ZN => n_679);
  g29640 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(0), B1 => n_462, B2 => snake_output21(0), ZN => n_678);
  g29641 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(3), B1 => n_539, B2 => n_1171, ZN => n_677);
  g29642 : ND4D0BWP7T port map(A1 => n_254, A2 => n_493, A3 => n_232, A4 => n_237, ZN => n_676);
  g29643 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(4), B1 => n_539, B2 => n_1172, ZN => n_675);
  g29644 : NR2D0BWP7T port map(A1 => n_610, A2 => n_438, ZN => n_700);
  g29645 : NR2D0BWP7T port map(A1 => n_619, A2 => corner_count(1), ZN => n_699);
  g29647 : INR2D0BWP7T port map(A1 => n_622, B1 => n_193, ZN => n_698);
  g29648 : NR2D0BWP7T port map(A1 => n_193, A2 => n_601, ZN => n_697);
  g29649 : NR3D0BWP7T port map(A1 => n_193, A2 => n_477, A3 => n_544, ZN => n_696);
  g29650 : NR2D0BWP7T port map(A1 => n_193, A2 => n_595, ZN => n_695);
  g29651 : NR2D0BWP7T port map(A1 => n_619, A2 => n_429, ZN => n_694);
  g29654 : NR2D0BWP7T port map(A1 => n_619, A2 => n_430, ZN => n_693);
  g29659 : OAI21D0BWP7T port map(A1 => n_541, A2 => n_217, B => n_195, ZN => n_765);
  g29660 : OAI21D0BWP7T port map(A1 => n_541, A2 => n_220, B => n_195, ZN => n_763);
  g29661 : AOI21D0BWP7T port map(A1 => n_565, A2 => n_212, B => n_194, ZN => n_762);
  g29662 : AOI21D0BWP7T port map(A1 => n_565, A2 => n_222, B => n_194, ZN => n_761);
  g29663 : AOI21D0BWP7T port map(A1 => n_564, A2 => n_222, B => n_194, ZN => n_759);
  g29665 : OAI21D0BWP7T port map(A1 => n_541, A2 => n_211, B => n_195, ZN => n_764);
  g29667 : IAO21D0BWP7T port map(A1 => n_566, A2 => n_220, B => n_194, ZN => n_757);
  g29669 : OAI21D0BWP7T port map(A1 => n_563, A2 => n_217, B => n_195, ZN => n_756);
  g29670 : AOI21D0BWP7T port map(A1 => n_565, A2 => n_218, B => n_194, ZN => n_758);
  g29672 : OAI21D0BWP7T port map(A1 => n_563, A2 => n_220, B => n_195, ZN => n_702);
  g29673 : AOI21D0BWP7T port map(A1 => n_564, A2 => n_212, B => n_194, ZN => n_760);
  g29674 : IOA21D0BWP7T port map(A1 => n_542, A2 => n_222, B => n_195, ZN => n_766);
  g29676 : NR2D0BWP7T port map(A1 => n_623, A2 => corner_count(0), ZN => n_692);
  g29677 : NR2D0BWP7T port map(A1 => n_623, A2 => n_146, ZN => n_691);
  g29678 : INR2D0BWP7T port map(A1 => n_425, B1 => n_619, ZN => n_690);
  g29679 : NR2D0BWP7T port map(A1 => n_619, A2 => n_428, ZN => n_689);
  g29680 : INR2D0BWP7T port map(A1 => n_622, B1 => n_478, ZN => n_688);
  g29681 : AN3D0BWP7T port map(A1 => n_477, A2 => n_544, A3 => n_420, Z => n_687);
  g29682 : NR3D0BWP7T port map(A1 => n_524, A2 => n_478, A3 => n_545, ZN => n_685);
  g29683 : AOI22D0BWP7T port map(A1 => n_546, A2 => snake_output17(5), B1 => n_462, B2 => snake_output22(5), ZN => n_672);
  g29684 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(0), B1 => n_496, B2 => snake_output1(0), ZN => n_671);
  g29685 : AOI22D0BWP7T port map(A1 => n_552, A2 => n_1120, B1 => n_418, B2 => snake_output14(0), ZN => n_670);
  g29686 : AOI22D0BWP7T port map(A1 => n_514, A2 => snake_output12(0), B1 => n_550, B2 => snake_output13(0), ZN => n_669);
  g29687 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(0), B1 => n_462, B2 => n_1066, ZN => n_668);
  g29688 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output10(0), B1 => n_514, B2 => snake_output11(0), ZN => n_667);
  g29689 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(1), B1 => n_462, B2 => snake_output21(1), ZN => n_666);
  g29690 : AOI22D0BWP7T port map(A1 => n_553, A2 => n_1049, B1 => n_559, B2 => snake_output16(1), ZN => n_665);
  g29691 : AOI22D0BWP7T port map(A1 => n_543, A2 => snake_output24(5), B1 => n_475, B2 => snake_output16(5), ZN => n_664);
  g29692 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(1), B1 => n_496, B2 => snake_output1(1), ZN => n_663);
  g29693 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output14(5), B1 => n_418, B2 => snake_output15(5), ZN => n_662);
  g29694 : AOI22D0BWP7T port map(A1 => n_552, A2 => n_1121, B1 => n_418, B2 => n_1103, ZN => n_661);
  g29695 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output12(5), B1 => n_514, B2 => snake_output13(5), ZN => n_660);
  g29696 : AOI22D0BWP7T port map(A1 => n_514, A2 => n_1115, B1 => n_550, B2 => n_1109, ZN => n_659);
  g29697 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(1), B1 => n_462, B2 => n_1067, ZN => n_658);
  g29698 : AOI22D0BWP7T port map(A1 => n_552, A2 => n_1127, B1 => n_514, B2 => snake_output11(1), ZN => n_657);
  g29699 : AOI22D0BWP7T port map(A1 => n_510, A2 => n_1181, B1 => n_532, B2 => snake_output5(1), ZN => n_656);
  g29700 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(2), B1 => n_462, B2 => snake_output21(2), ZN => n_655);
  g29701 : AOI22D0BWP7T port map(A1 => n_553, A2 => n_1050, B1 => n_559, B2 => snake_output16(2), ZN => n_654);
  g29702 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(2), B1 => n_496, B2 => snake_output1(2), ZN => n_653);
  g29703 : AOI22D0BWP7T port map(A1 => n_555, A2 => n_1185, B1 => n_507, B2 => snake_output0(5), ZN => n_652);
  g29704 : AOI22D0BWP7T port map(A1 => n_552, A2 => n_1122, B1 => n_418, B2 => snake_output14(2), ZN => n_651);
  g29705 : AOI22D0BWP7T port map(A1 => n_514, A2 => n_1116, B1 => n_550, B2 => snake_output13(2), ZN => n_650);
  g29706 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(2), B1 => n_462, B2 => n_1068, ZN => n_649);
  g29707 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output12(2), B1 => n_418, B2 => n_1110, ZN => n_648);
  g29708 : AOI22D0BWP7T port map(A1 => n_510, A2 => n_1182, B1 => n_532, B2 => snake_output5(2), ZN => n_647);
  g29709 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(3), B1 => n_462, B2 => snake_output21(3), ZN => n_646);
  g29710 : AOI22D0BWP7T port map(A1 => n_553, A2 => n_1051, B1 => n_559, B2 => snake_output16(3), ZN => n_645);
  g29711 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(3), B1 => n_496, B2 => snake_output1(3), ZN => n_644);
  g29712 : AOI22D0BWP7T port map(A1 => n_514, A2 => n_1117, B1 => n_550, B2 => snake_output13(3), ZN => n_643);
  g29713 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(3), B1 => n_462, B2 => n_1069, ZN => n_642);
  g29714 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output12(3), B1 => n_418, B2 => n_1111, ZN => n_641);
  g29715 : AOI22D0BWP7T port map(A1 => n_500, A2 => n_1165, B1 => n_532, B2 => snake_output5(3), ZN => n_640);
  g29716 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(4), B1 => n_462, B2 => snake_output21(4), ZN => n_639);
  g29717 : AOI22D0BWP7T port map(A1 => n_553, A2 => n_1052, B1 => n_559, B2 => snake_output16(4), ZN => n_638);
  g29718 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(4), B1 => n_496, B2 => snake_output1(4), ZN => n_637);
  g29719 : AOI22D0BWP7T port map(A1 => n_552, A2 => n_1124, B1 => n_418, B2 => snake_output14(4), ZN => n_636);
  g29720 : AOI22D0BWP7T port map(A1 => n_514, A2 => n_1118, B1 => n_550, B2 => snake_output13(4), ZN => n_635);
  g29721 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(4), B1 => n_462, B2 => n_1070, ZN => n_634);
  g29722 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output12(4), B1 => n_418, B2 => n_1112, ZN => n_633);
  g29723 : AOI22D0BWP7T port map(A1 => n_552, A2 => n_1123, B1 => n_418, B2 => snake_output14(3), ZN => n_632);
  g29724 : AOI22D0BWP7T port map(A1 => n_510, A2 => n_1184, B1 => n_532, B2 => snake_output5(4), ZN => n_631);
  g29725 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output6(5), B1 => n_532, B2 => snake_output7(5), ZN => n_630);
  g29726 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(0), B1 => n_550, B2 => n_1114, ZN => n_629);
  g29727 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(1), B1 => n_550, B2 => snake_output12(1), ZN => n_628);
  g29728 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(2), B1 => n_552, B2 => snake_output10(2), ZN => n_627);
  g29729 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(3), B1 => n_552, B2 => snake_output10(3), ZN => n_626);
  g29730 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(4), B1 => n_552, B2 => snake_output10(4), ZN => n_625);
  g29731 : AOI22D0BWP7T port map(A1 => n_553, A2 => n_1048, B1 => n_559, B2 => snake_output16(0), ZN => n_624);
  g29733 : CKND1BWP7T port map(I => n_602, ZN => n_601);
  g29734 : OAI31D0BWP7T port map(A1 => N(0), A2 => n_230, A3 => n_423, B => n_232, ZN => n_600);
  g29735 : AOI31D0BWP7T port map(A1 => n_485, A2 => N(0), A3 => n_1185, B => n_489, ZN => n_599);
  g29736 : ND2D0BWP7T port map(A1 => n_536, A2 => n_228, ZN => n_623);
  g29737 : NR2D0BWP7T port map(A1 => n_523, A2 => n_545, ZN => n_622);
  g29738 : AN2D1BWP7T port map(A1 => n_478, A2 => n_545, Z => n_621);
  g29739 : INR2D0BWP7T port map(A1 => n_546, B1 => n_193, ZN => n_620);
  g29740 : ND2D0BWP7T port map(A1 => n_535, A2 => n_463, ZN => n_619);
  g29741 : INR2D0BWP7T port map(A1 => n_554, B1 => n_193, ZN => n_618);
  g29742 : INR2D0BWP7T port map(A1 => n_554, B1 => n_478, ZN => n_617);
  g29743 : NR2D0BWP7T port map(A1 => n_193, A2 => n_549, ZN => n_616);
  g29744 : NR2D0BWP7T port map(A1 => n_193, A2 => n_531, ZN => n_615);
  g29745 : INR2D0BWP7T port map(A1 => n_555, B1 => n_193, ZN => n_614);
  g29746 : NR2D0BWP7T port map(A1 => n_193, A2 => n_551, ZN => n_613);
  g29747 : NR2D0BWP7T port map(A1 => n_193, A2 => n_533, ZN => n_612);
  g29748 : AOI211D0BWP7T port map(A1 => n_485, A2 => N(4), B => n_464, C => n_508, ZN => n_611);
  g29750 : ND2D0BWP7T port map(A1 => n_529, A2 => n_1698, ZN => n_610);
  g29751 : INR2D0BWP7T port map(A1 => n_425, B1 => n_535, ZN => n_609);
  g29753 : NR2D0BWP7T port map(A1 => n_535, A2 => n_428, ZN => n_608);
  g29755 : NR2D0BWP7T port map(A1 => n_535, A2 => n_435, ZN => n_607);
  g29758 : NR2D0BWP7T port map(A1 => n_535, A2 => n_436, ZN => n_606);
  g29759 : NR2D0BWP7T port map(A1 => n_535, A2 => n_430, ZN => n_605);
  g29760 : NR2D0BWP7T port map(A1 => n_535, A2 => n_463, ZN => n_604);
  g29762 : NR3D0BWP7T port map(A1 => n_429, A2 => n_536, A3 => n_463, ZN => n_603);
  g29763 : OAI21D0BWP7T port map(A1 => n_522, A2 => n_1700, B => n_195, ZN => n_674);
  g29764 : NR4D0BWP7T port map(A1 => n_477, A2 => n_466, A3 => n_421, A4 => N(0), ZN => n_602);
  g29765 : INVD0BWP7T port map(I => n_596, ZN => n_595);
  g29766 : AOI22D0BWP7T port map(A1 => n_498, A2 => n_1177, B1 => n_510, B2 => n_1183, ZN => n_594);
  g29767 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(1), B1 => n_519, B2 => n_1121, ZN => n_593);
  g29768 : AOI22D0BWP7T port map(A1 => n_520, A2 => n_1115, B1 => n_505, B2 => snake_output13(1), ZN => n_592);
  g29769 : AOI22D0BWP7T port map(A1 => n_504, A2 => n_1128, B1 => n_519, B2 => n_1122, ZN => n_591);
  g29770 : AOI22D0BWP7T port map(A1 => n_512, A2 => n_1126, B1 => n_475, B2 => n_1096, ZN => n_590);
  g29771 : AOI22D0BWP7T port map(A1 => n_506, A2 => n_1090, B1 => n_502, B2 => n_1072, ZN => n_589);
  g29772 : AOI22D0BWP7T port map(A1 => n_500, A2 => n_1162, B1 => n_496, B2 => snake_output0(0), ZN => n_588);
  g29773 : AOI22D0BWP7T port map(A1 => n_512, A2 => n_1127, B1 => n_475, B2 => n_1097, ZN => n_587);
  g29774 : AOI22D0BWP7T port map(A1 => n_506, A2 => n_1091, B1 => n_502, B2 => n_1073, ZN => n_586);
  g29775 : AOI22D0BWP7T port map(A1 => n_500, A2 => n_1163, B1 => n_496, B2 => snake_output0(1), ZN => n_585);
  g29776 : AOI22D0BWP7T port map(A1 => n_498, A2 => n_1167, B1 => n_510, B2 => snake_output3(5), ZN => n_584);
  g29777 : AOI22D0BWP7T port map(A1 => n_512, A2 => n_1128, B1 => n_475, B2 => n_1098, ZN => n_583);
  g29778 : AOI22D0BWP7T port map(A1 => n_506, A2 => n_1092, B1 => n_502, B2 => n_1074, ZN => n_582);
  g29779 : AOI22D0BWP7T port map(A1 => n_500, A2 => n_1164, B1 => n_496, B2 => snake_output0(2), ZN => n_581);
  g29780 : AOI22D0BWP7T port map(A1 => n_512, A2 => n_1129, B1 => n_475, B2 => n_1099, ZN => n_580);
  g29781 : AOI22D0BWP7T port map(A1 => n_506, A2 => n_1093, B1 => n_502, B2 => n_1075, ZN => n_579);
  g29782 : AOI22D0BWP7T port map(A1 => n_520, A2 => n_1116, B1 => n_505, B2 => n_1110, ZN => n_578);
  g29783 : AOI22D0BWP7T port map(A1 => n_512, A2 => n_1130, B1 => n_475, B2 => n_1100, ZN => n_577);
  g29784 : AOI22D0BWP7T port map(A1 => n_506, A2 => n_1094, B1 => n_502, B2 => n_1076, ZN => n_576);
  g29785 : AOI22D0BWP7T port map(A1 => n_500, A2 => n_1166, B1 => n_496, B2 => snake_output0(4), ZN => n_575);
  g29786 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(5), B1 => n_519, B2 => n_1125, ZN => n_574);
  g29787 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(5), B1 => n_505, B2 => snake_output13(5), ZN => n_573);
  g29788 : AOI22D0BWP7T port map(A1 => n_520, A2 => n_1118, B1 => n_505, B2 => n_1112, ZN => n_572);
  g29789 : AOI22D0BWP7T port map(A1 => n_504, A2 => n_1130, B1 => n_519, B2 => n_1124, ZN => n_571);
  g29790 : AOI22D0BWP7T port map(A1 => n_520, A2 => n_1117, B1 => n_505, B2 => n_1111, ZN => n_570);
  g29791 : AOI22D0BWP7T port map(A1 => n_504, A2 => n_1129, B1 => n_519, B2 => n_1123, ZN => n_569);
  g29792 : AOI22D0BWP7T port map(A1 => n_504, A2 => n_1126, B1 => n_519, B2 => n_1120, ZN => n_568);
  g29793 : AOI22D0BWP7T port map(A1 => n_520, A2 => n_1114, B1 => n_505, B2 => n_1108, ZN => n_567);
  g29794 : AO21D0BWP7T port map(A1 => n_192, A2 => n_507, B => n_1737, Z => n_597);
  g29795 : IAO21D0BWP7T port map(A1 => n_522, A2 => n_150, B => n_194, ZN => n_673);
  g29797 : INR4D0BWP7T port map(A1 => n_466, B1 => N(0), B2 => n_421, B3 => n_477, ZN => n_596);
  g29798 : CKND1BWP7T port map(I => n_565, ZN => n_566);
  g29799 : CKND1BWP7T port map(I => n_564, ZN => n_563);
  g29800 : CKND1BWP7T port map(I => n_552, ZN => n_551);
  g29801 : CKND1BWP7T port map(I => n_550, ZN => n_549);
  g29803 : NR2D0BWP7T port map(A1 => n_492, A2 => n_230, ZN => n_547);
  g29804 : NR2D0BWP7T port map(A1 => n_525, A2 => n_1701, ZN => n_565);
  g29805 : NR2D0BWP7T port map(A1 => n_525, A2 => n_156, ZN => n_564);
  g29806 : NR2D0BWP7T port map(A1 => n_523, A2 => n_479, ZN => n_562);
  g29807 : NR2D0BWP7T port map(A1 => n_193, A2 => n_499, ZN => n_561);
  g29808 : NR2D0BWP7T port map(A1 => n_193, A2 => n_501, ZN => n_560);
  g29809 : AN2D1BWP7T port map(A1 => n_503, A2 => N(4), Z => n_559);
  g29810 : NR2D0BWP7T port map(A1 => n_193, A2 => n_513, ZN => n_558);
  g29811 : NR2D0BWP7T port map(A1 => n_193, A2 => n_511, ZN => n_557);
  g29812 : INR2D0BWP7T port map(A1 => n_515, B1 => n_193, ZN => n_556);
  g29813 : AN2D1BWP7T port map(A1 => n_503, A2 => n_477, Z => n_555);
  g29814 : NR2D0BWP7T port map(A1 => n_521, A2 => n_224, ZN => n_554);
  g29815 : NR2D0BWP7T port map(A1 => n_524, A2 => n_479, ZN => n_553);
  g29816 : INR2D0BWP7T port map(A1 => n_226, B1 => n_521, ZN => n_552);
  g29817 : NR2D0BWP7T port map(A1 => n_521, A2 => n_221, ZN => n_550);
  g29818 : INVD0BWP7T port map(I => n_544, ZN => n_543);
  g29819 : CKND1BWP7T port map(I => n_541, ZN => n_542);
  g29820 : INVD1BWP7T port map(I => n_536, ZN => n_535);
  g29821 : CKND1BWP7T port map(I => n_534, ZN => n_533);
  g29822 : INVD1BWP7T port map(I => n_531, ZN => n_532);
  g29823 : INR4D0BWP7T port map(A1 => n_452, B1 => n_1734, B2 => n_1739, B3 => n_1737, ZN => n_530);
  g29824 : NR4D0BWP7T port map(A1 => n_469, A2 => n_1695, A3 => n_1696, A4 => n_1697, ZN => n_529);
  g29825 : INR4D0BWP7T port map(A1 => n_449, B1 => corner_count(31), B2 => corner_count(30), B3 => corner_count(29), ZN => n_528);
  g29826 : AOI22D0BWP7T port map(A1 => n_475, A2 => n_1102, B1 => n_418, B2 => n_1108, ZN => n_527);
  g29827 : AOI31D0BWP7T port map(A1 => n_214, A2 => N(3), A3 => n_1047, B => n_491, ZN => n_526);
  g29828 : AN3D0BWP7T port map(A1 => n_476, A2 => n_468, A3 => n_466, Z => n_546);
  g29829 : OAI21D0BWP7T port map(A1 => n_484, A2 => n_149, B => n_424, ZN => n_545);
  g29830 : AOI21D0BWP7T port map(A1 => n_488, A2 => N(3), B => n_418, ZN => n_544);
  g29831 : IND3D0BWP7T port map(A1 => n_1699, B1 => n_1701, B2 => n_481, ZN => n_541);
  g29832 : NR2D0BWP7T port map(A1 => n_193, A2 => n_497, ZN => n_540);
  g29833 : NR2D0BWP7T port map(A1 => n_193, A2 => n_509, ZN => n_539);
  g29834 : NR3D0BWP7T port map(A1 => n_193, A2 => n_474, A3 => n_477, ZN => n_538);
  g29835 : NR2D0BWP7T port map(A1 => n_193, A2 => n_495, ZN => n_537);
  g29836 : IAO21D0BWP7T port map(A1 => n_482, A2 => n_434, B => n_194, ZN => n_598);
  g29837 : CKXOR2D0BWP7T port map(A1 => corner_count(4), A2 => n_419, Z => n_536);
  g29838 : NR3D0BWP7T port map(A1 => n_467, A2 => n_466, A3 => n_147, ZN => n_534);
  g29839 : ND3D0BWP7T port map(A1 => n_426, A2 => n_147, A3 => N(3), ZN => n_531);
  g29840 : CKND1BWP7T port map(I => n_514, ZN => n_513);
  g29841 : CKND1BWP7T port map(I => n_512, ZN => n_511);
  g29842 : CKND1BWP7T port map(I => n_510, ZN => n_509);
  g29843 : NR2D0BWP7T port map(A1 => n_485, A2 => N(4), ZN => n_508);
  g29844 : ND2D0BWP7T port map(A1 => n_481, A2 => n_1699, ZN => n_525);
  g29845 : OR2D0BWP7T port map(A1 => n_467, A2 => n_486, Z => n_524);
  g29846 : ND2D0BWP7T port map(A1 => n_468, A2 => n_487, ZN => n_523);
  g29847 : IND2D0BWP7T port map(A1 => n_438, B1 => n_481, ZN => n_522);
  g29848 : IND2D0BWP7T port map(A1 => n_464, B1 => N(0), ZN => n_521);
  g29849 : INR2D0BWP7T port map(A1 => n_425, B1 => n_463, ZN => n_520);
  g29850 : NR2D0BWP7T port map(A1 => n_435, A2 => n_463, ZN => n_519);
  g29851 : INR2D0BWP7T port map(A1 => n_419, B1 => n_146, ZN => n_518);
  g29852 : INR2D0BWP7T port map(A1 => n_419, B1 => corner_count(0), ZN => n_517);
  g29853 : NR2D0BWP7T port map(A1 => n_428, A2 => n_463, ZN => n_516);
  g29854 : NR2D0BWP7T port map(A1 => n_487, A2 => n_439, ZN => n_515);
  g29855 : INR2D0BWP7T port map(A1 => n_420, B1 => n_464, ZN => n_514);
  g29856 : NR2D0BWP7T port map(A1 => n_464, A2 => n_433, ZN => n_512);
  g29857 : NR2D0BWP7T port map(A1 => n_478, A2 => n_437, ZN => n_510);
  g29858 : INVD1BWP7T port map(I => n_501, ZN => n_502);
  g29859 : CKND1BWP7T port map(I => n_500, ZN => n_499);
  g29860 : CKND1BWP7T port map(I => n_498, ZN => n_497);
  g29861 : CKND1BWP7T port map(I => n_496, ZN => n_495);
  g29862 : AOI33D0BWP7T port map(A1 => n_432, A2 => n_214, A3 => n_1071, B1 => n_420, B2 => n_223, B3 => n_1107, ZN => n_494);
  g29863 : MAOI22D0BWP7T port map(A1 => n_1572, A2 => n_448, B1 => n_154, B2 => send_corner_flag, ZN => n_493);
  g29864 : AOI31D0BWP7T port map(A1 => n_420, A2 => n_149, A3 => n_1155, B => n_457, ZN => n_492);
  g29865 : NR3D0BWP7T port map(A1 => n_460, A2 => n_224, A3 => N(0), ZN => n_491);
  g29866 : AOI22D0BWP7T port map(A1 => n_442, A2 => n_427, B1 => n_458, B2 => n_1119, ZN => n_490);
  g29867 : OAI32D0BWP7T port map(A1 => n_153, A2 => n_215, A3 => n_239, B1 => n_144, B2 => n_437, ZN => n_489);
  g29868 : NR2D0BWP7T port map(A1 => n_474, A2 => n_476, ZN => n_507);
  g29869 : NR2D0BWP7T port map(A1 => n_479, A2 => n_441, ZN => n_506);
  g29870 : NR2D0BWP7T port map(A1 => n_430, A2 => n_463, ZN => n_505);
  g29871 : NR2D0BWP7T port map(A1 => n_436, A2 => n_463, ZN => n_504);
  g29872 : AN3D0BWP7T port map(A1 => n_464, A2 => n_468, A3 => n_221, Z => n_503);
  g29873 : ND2D0BWP7T port map(A1 => n_476, A2 => n_420, ZN => n_501);
  g29874 : NR3D0BWP7T port map(A1 => n_478, A2 => n_421, A3 => n_431, ZN => n_500);
  g29875 : NR3D0BWP7T port map(A1 => n_476, A2 => n_422, A3 => n_431, ZN => n_498);
  g29876 : NR2D0BWP7T port map(A1 => n_478, A2 => n_441, ZN => n_496);
  g29877 : CKND1BWP7T port map(I => n_426, ZN => n_488);
  g29879 : INVD0BWP7T port map(I => n_486, ZN => n_487);
  g29880 : CKND1BWP7T port map(I => n_423, ZN => n_485);
  g29881 : HA1D0BWP7T port map(A => n_148, B => n_210, CO => n_484, S => n_486);
  g29902 : CKND1BWP7T port map(I => n_481, ZN => n_482);
  g29903 : INVD1BWP7T port map(I => n_479, ZN => n_478);
  g29904 : INVD1BWP7T port map(I => n_477, ZN => n_476);
  g29905 : CKND1BWP7T port map(I => n_475, ZN => n_474);
  g29913 : AOI22D0BWP7T port map(A1 => n_418, A2 => n_1095, B1 => n_420, B2 => n_1059, ZN => n_473);
  g29918 : MAOI22D0BWP7T port map(A1 => n_427, A2 => n_1101, B1 => n_440, B2 => n_145, ZN => n_472);
  g29920 : AOI222D0BWP7T port map(A1 => n_219, A2 => n_1089, B1 => n_226, B2 => snake_output21(5), C1 => n_225, C2 => n_1077, ZN => n_471);
  g29921 : NR2D0BWP7T port map(A1 => n_469, A2 => n_1582, ZN => n_481);
  g29922 : NR2D0BWP7T port map(A1 => n_193, A2 => n_461, ZN => n_480);
  g29923 : MAOI22D0BWP7T port map(A1 => n_424, A2 => N(4), B1 => n_424, B2 => N(4), ZN => n_479);
  g29925 : AOI22D0BWP7T port map(A1 => n_418, A2 => n_147, B1 => n_417, B2 => N(4), ZN => n_477);
  g29926 : NR2D0BWP7T port map(A1 => n_467, A2 => n_215, ZN => n_475);
  g29956 : CKND1BWP7T port map(I => n_462, ZN => n_461);
  g29957 : AOI22D0BWP7T port map(A1 => n_214, A2 => n_1083, B1 => n_223, B2 => n_1131, ZN => n_460);
  g29958 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(4), B1 => n_207, B2 => snake_output0(4), ZN => n_459);
  g29959 : INR2D0BWP7T port map(A1 => n_223, B1 => n_433, ZN => n_458);
  g29960 : NR2D0BWP7T port map(A1 => n_431, A2 => n_238, ZN => n_457);
  g29961 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(3), B1 => n_207, B2 => snake_output0(3), ZN => n_456);
  g29962 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(1), B1 => n_207, B2 => snake_output0(1), ZN => n_455);
  g29963 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(0), B1 => n_207, B2 => snake_output0(0), ZN => n_454);
  g29964 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(2), B1 => n_1737, B2 => head(7), ZN => n_453);
  g29965 : NR4D0BWP7T port map(A1 => n_1579, A2 => n_1735, A3 => n_1736, A4 => n_1738, ZN => n_452);
  g29966 : AO221D0BWP7T port map(A1 => n_1703, A2 => n_146, B1 => n_1704, B2 => new_corner_count(0), C => n_1739, Z => n_451);
  g29967 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(4), B1 => n_207, B2 => head(9), ZN => n_450);
  g29968 : NR4D0BWP7T port map(A1 => corner_count(16), A2 => corner_count(15), A3 => corner_count(14), A4 => corner_count(13), ZN => n_449);
  g29969 : AO211D0BWP7T port map(A1 => n_1273, A2 => n_1742, B => n_1575, C => new_head_flag, Z => n_448);
  g29970 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(3), B1 => n_207, B2 => head(8), ZN => n_447);
  g29971 : IIND4D0BWP7T port map(A1 => n_1573, A2 => n_1574, B1 => n_1572, B2 => n_1585, ZN => n_446);
  g29972 : AOI22D0BWP7T port map(A1 => n_207, A2 => head(7), B1 => n_1737, B2 => head(2), ZN => n_445);
  g29973 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(1), B1 => n_207, B2 => head(6), ZN => n_444);
  g29974 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(0), B1 => n_207, B2 => head(5), ZN => n_443);
  g29975 : AO22D0BWP7T port map(A1 => n_219, A2 => snake_output9(5), B1 => snake_output11(5), B2 => n_225, Z => n_442);
  g29976 : OAI211D0BWP7T port map(A1 => n_1670, A2 => n_1703, B => n_1580, C => n_187, ZN => n_469);
  g29978 : NR2D0BWP7T port map(A1 => n_422, A2 => N(0), ZN => n_468);
  g29979 : ND2D0BWP7T port map(A1 => n_421, A2 => N(0), ZN => n_467);
  g29981 : AOI21D0BWP7T port map(A1 => n_216, A2 => N(2), B => n_426, ZN => n_466);
  g29982 : NR2D0BWP7T port map(A1 => n_193, A2 => n_417, ZN => n_465);
  g29983 : OA21D0BWP7T port map(A1 => n_219, A2 => n_149, B => n_423, Z => n_464);
  g29984 : AOI21D0BWP7T port map(A1 => n_229, A2 => corner_count(3), B => n_419, ZN => n_463);
  g29985 : NR2D0BWP7T port map(A1 => n_439, A2 => n_148, ZN => n_462);
  g29986 : NR4D0BWP7T port map(A1 => n_1739, A2 => n_1734, A3 => n_1662, A4 => n_1736, ZN => n_483);
  g29987 : INVD0BWP7T port map(I => n_433, ZN => n_432);
  g29988 : INVD1BWP7T port map(I => n_422, ZN => n_421);
  g29989 : INVD1BWP7T port map(I => n_418, ZN => n_417);
  g29995 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift9(1), B => n_201, ZN => n_416);
  g29996 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift8(5), B => n_197, ZN => n_415);
  g29997 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift8(3), B => n_198, ZN => n_414);
  g29998 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift5(3), B => n_198, ZN => n_413);
  g29999 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift8(1), B => n_201, ZN => n_412);
  g30000 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift7(5), B => n_197, ZN => n_411);
  g30001 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(5), B => n_197, ZN => n_410);
  g30002 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift7(4), B => n_196, ZN => n_409);
  g30003 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift7(3), B => n_198, ZN => n_408);
  g30004 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift16(0), B => n_199, ZN => n_407);
  g30005 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift6(0), B => n_199, ZN => n_406);
  g30006 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift7(1), B => n_201, ZN => n_405);
  g30007 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift6(4), B => n_196, ZN => n_404);
  g30008 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift6(3), B => n_198, ZN => n_403);
  g30009 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift6(2), B => n_200, ZN => n_402);
  g30010 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift4(1), B => n_201, ZN => n_401);
  g30011 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift8(2), B => n_200, ZN => n_400);
  g30012 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift6(1), B => n_201, ZN => n_399);
  g30013 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift4(2), B => n_200, ZN => n_398);
  g30014 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift8(0), B => n_199, ZN => n_397);
  g30015 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(0), B => n_199, ZN => n_396);
  g30016 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift4(4), B => n_196, ZN => n_395);
  g30017 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift4(0), B => n_199, ZN => n_394);
  g30018 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(1), B => n_201, ZN => n_393);
  g30019 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift19(0), B => n_199, ZN => n_392);
  g30020 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift19(1), B => n_201, ZN => n_391);
  g30021 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift19(2), B => n_200, ZN => n_390);
  g30022 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift19(3), B => n_198, ZN => n_389);
  g30023 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(2), B => n_200, ZN => n_388);
  g30024 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift19(4), B => n_196, ZN => n_387);
  g30025 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(3), B => n_198, ZN => n_386);
  g30026 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift19(5), B => n_197, ZN => n_385);
  g30027 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift20(0), B => n_199, ZN => n_384);
  g30028 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift20(1), B => n_201, ZN => n_383);
  g30029 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift20(2), B => n_200, ZN => n_382);
  g30030 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(4), B => n_196, ZN => n_381);
  g30031 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift20(3), B => n_198, ZN => n_380);
  g30032 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift20(4), B => n_196, ZN => n_379);
  g30033 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift20(5), B => n_197, ZN => n_378);
  g30034 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift21(0), B => n_199, ZN => n_377);
  g30035 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(0), B => n_199, ZN => n_376);
  g30036 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift4(5), B => n_197, ZN => n_375);
  g30037 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(5), B => n_197, ZN => n_374);
  g30038 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift21(1), B => n_201, ZN => n_373);
  g30039 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift21(2), B => n_200, ZN => n_372);
  g30040 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift21(3), B => n_198, ZN => n_371);
  g30041 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(2), B => n_200, ZN => n_370);
  g30042 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift22(0), B => n_199, ZN => n_369);
  g30043 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift22(1), B => n_201, ZN => n_368);
  g30044 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(3), B => n_198, ZN => n_367);
  g30045 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift22(2), B => n_200, ZN => n_366);
  g30046 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift22(4), B => n_196, ZN => n_365);
  g30047 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift22(5), B => n_197, ZN => n_364);
  g30048 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(4), B => n_196, ZN => n_363);
  g30049 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift23(0), B => n_199, ZN => n_362);
  g30050 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift23(1), B => n_201, ZN => n_361);
  g30051 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift8(4), B => n_196, ZN => n_360);
  g30052 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift23(4), B => n_196, ZN => n_359);
  g30053 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift23(3), B => n_198, ZN => n_358);
  g30054 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift23(5), B => n_197, ZN => n_357);
  g30055 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(5), B => n_197, ZN => n_356);
  g30056 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(2), B => n_200, ZN => n_355);
  g30057 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift5(4), B => n_196, ZN => n_354);
  g30058 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(1), B => n_201, ZN => n_353);
  g30059 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(4), B => n_196, ZN => n_352);
  g30060 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift23(2), B => n_200, ZN => n_351);
  g30061 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(5), B => n_197, ZN => n_350);
  g30062 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(0), B => n_199, ZN => n_349);
  g30063 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(1), B => n_201, ZN => n_348);
  g30064 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift21(5), B => n_197, ZN => n_347);
  g30065 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift21(4), B => n_196, ZN => n_346);
  g30066 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(2), B => n_200, ZN => n_345);
  g30067 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(3), B => n_198, ZN => n_344);
  g30068 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(4), B => n_196, ZN => n_343);
  g30069 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift7(0), B => n_199, ZN => n_342);
  g30070 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift22(3), B => n_198, ZN => n_341);
  g30071 : OR2D0BWP7T port map(A1 => n_210, A2 => n_215, Z => n_441);
  g30072 : ND2D0BWP7T port map(A1 => n_214, A2 => N(0), ZN => n_440);
  g30073 : IND2D0BWP7T port map(A1 => n_210, B1 => N(4), ZN => n_439);
  g30074 : ND2D0BWP7T port map(A1 => n_235, A2 => n_146, ZN => n_438);
  g30075 : IND2D0BWP7T port map(A1 => n_216, B1 => n_234, ZN => n_437);
  g30076 : IND2D0BWP7T port map(A1 => corner_count(1), B1 => n_231, ZN => n_436);
  g30077 : IND2D0BWP7T port map(A1 => corner_count(1), B1 => n_227, ZN => n_435);
  g30078 : ND2D0BWP7T port map(A1 => n_235, A2 => n_218, ZN => n_434);
  g30079 : ND2D0BWP7T port map(A1 => n_226, A2 => n_152, ZN => n_433);
  g30080 : ND2D0BWP7T port map(A1 => n_234, A2 => N(0), ZN => n_431);
  g30081 : IND2D0BWP7T port map(A1 => n_233, B1 => corner_count(0), ZN => n_430);
  g30082 : ND2D0BWP7T port map(A1 => n_231, A2 => corner_count(1), ZN => n_429);
  g30083 : ND2D0BWP7T port map(A1 => n_227, A2 => corner_count(1), ZN => n_428);
  g30084 : AN2D1BWP7T port map(A1 => n_223, A2 => N(0), Z => n_427);
  g30085 : NR2D0BWP7T port map(A1 => n_216, A2 => N(2), ZN => n_426);
  g30086 : NR2D0BWP7T port map(A1 => n_233, A2 => corner_count(0), ZN => n_425);
  g30087 : IND2D0BWP7T port map(A1 => n_215, B1 => n_210, ZN => n_424);
  g30088 : ND2D0BWP7T port map(A1 => n_219, A2 => n_149, ZN => n_423);
  g30089 : ND2D0BWP7T port map(A1 => n_210, A2 => n_216, ZN => n_422);
  g30090 : NR2D0BWP7T port map(A1 => n_221, A2 => N(0), ZN => n_420);
  g30091 : NR2D0BWP7T port map(A1 => n_229, A2 => corner_count(3), ZN => n_419);
  g30092 : NR2D0BWP7T port map(A1 => n_215, A2 => n_216, ZN => n_418);
  g30093 : NR2D0BWP7T port map(A1 => n_194, A2 => n_1703, ZN => n_470);
  g30094 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift9(2), B => n_200, ZN => n_340);
  g30095 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift9(3), B => n_198, ZN => n_339);
  g30096 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift9(4), B => n_196, ZN => n_338);
  g30097 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift9(5), B => n_197, ZN => n_337);
  g30098 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift10(0), B => n_199, ZN => n_336);
  g30099 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift4(3), B => n_198, ZN => n_335);
  g30100 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift10(1), B => n_201, ZN => n_334);
  g30101 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift10(2), B => n_200, ZN => n_333);
  g30102 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift10(3), B => n_198, ZN => n_332);
  g30103 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift10(4), B => n_196, ZN => n_331);
  g30104 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift10(5), B => n_197, ZN => n_330);
  g30105 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift11(0), B => n_199, ZN => n_329);
  g30106 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift9(0), B => n_199, ZN => n_328);
  g30107 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift11(1), B => n_201, ZN => n_327);
  g30108 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift11(2), B => n_200, ZN => n_326);
  g30109 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift11(3), B => n_198, ZN => n_325);
  g30110 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift11(4), B => n_196, ZN => n_324);
  g30111 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift11(5), B => n_197, ZN => n_323);
  g30112 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift12(0), B => n_199, ZN => n_322);
  g30113 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift5(0), B => n_199, ZN => n_321);
  g30114 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift12(1), B => n_201, ZN => n_320);
  g30115 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift7(2), B => n_200, ZN => n_319);
  g30116 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift12(2), B => n_200, ZN => n_318);
  g30117 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift12(3), B => n_198, ZN => n_317);
  g30118 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift12(4), B => n_196, ZN => n_316);
  g30119 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift12(5), B => n_197, ZN => n_315);
  g30120 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift13(0), B => n_199, ZN => n_314);
  g30121 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift13(1), B => n_201, ZN => n_313);
  g30122 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift13(2), B => n_200, ZN => n_312);
  g30123 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift13(3), B => n_198, ZN => n_311);
  g30124 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift13(4), B => n_196, ZN => n_310);
  g30125 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift13(5), B => n_197, ZN => n_309);
  g30126 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift6(5), B => n_197, ZN => n_308);
  g30127 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift14(0), B => n_199, ZN => n_307);
  g30128 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift14(1), B => n_201, ZN => n_306);
  g30129 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift14(2), B => n_200, ZN => n_305);
  g30130 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift14(3), B => n_198, ZN => n_304);
  g30131 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift14(4), B => n_196, ZN => n_303);
  g30132 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift14(5), B => n_197, ZN => n_302);
  g30133 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift15(0), B => n_199, ZN => n_301);
  g30134 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift15(1), B => n_201, ZN => n_300);
  g30135 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift15(2), B => n_200, ZN => n_299);
  g30136 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(1), B => n_201, ZN => n_298);
  g30137 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift15(3), B => n_198, ZN => n_297);
  g30138 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift15(4), B => n_196, ZN => n_296);
  g30139 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift15(5), B => n_197, ZN => n_295);
  g30140 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(3), B => n_198, ZN => n_294);
  g30141 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift16(1), B => n_201, ZN => n_293);
  g30142 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift16(2), B => n_200, ZN => n_292);
  g30143 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift16(3), B => n_198, ZN => n_291);
  g30144 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift16(4), B => n_196, ZN => n_290);
  g30145 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift16(5), B => n_197, ZN => n_289);
  g30146 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift5(5), B => n_197, ZN => n_288);
  g30147 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift17(0), B => n_199, ZN => n_287);
  g30148 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift5(2), B => n_200, ZN => n_286);
  g30149 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift17(1), B => n_201, ZN => n_285);
  g30150 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift5(1), B => n_201, ZN => n_284);
  g30151 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift17(2), B => n_200, ZN => n_283);
  g30152 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift17(3), B => n_198, ZN => n_282);
  g30153 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift17(4), B => n_196, ZN => n_281);
  g30154 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift17(5), B => n_197, ZN => n_280);
  g30155 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(0), B => n_199, ZN => n_279);
  g30156 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift18(0), B => n_199, ZN => n_278);
  g30157 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift18(1), B => n_201, ZN => n_277);
  g30158 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift18(2), B => n_200, ZN => n_276);
  g30159 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift18(3), B => n_198, ZN => n_275);
  g30160 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift18(4), B => n_196, ZN => n_274);
  g30161 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift18(5), B => n_197, ZN => n_273);
  g30162 : AO22D0BWP7T port map(A1 => n_1693, A2 => n_1703, B1 => new_corner_count(9), B2 => n_1704, Z => n_272);
  g30163 : AO22D0BWP7T port map(A1 => n_1692, A2 => n_1703, B1 => new_corner_count(10), B2 => n_1704, Z => n_271);
  g30164 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1698, B1 => new_corner_count(4), B2 => n_1704, Z => n_270);
  g30165 : MOAI22D0BWP7T port map(A1 => n_151, A2 => n_150, B1 => n_1704, B2 => new_corner_count(2), ZN => n_269);
  g30166 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1699, B1 => new_corner_count(3), B2 => n_1704, Z => n_268);
  g30167 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1697, B1 => new_corner_count(5), B2 => n_1704, Z => n_267);
  g30168 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1696, B1 => new_corner_count(6), B2 => n_1704, Z => n_266);
  g30169 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1695, B1 => new_corner_count(7), B2 => n_1704, Z => n_265);
  g30170 : AO22D0BWP7T port map(A1 => n_1694, A2 => n_1703, B1 => new_corner_count(8), B2 => n_1704, Z => n_264);
  g30171 : AO22D0BWP7T port map(A1 => n_1680, A2 => n_1703, B1 => new_corner_count(22), B2 => n_1704, Z => n_263);
  g30172 : AO22D0BWP7T port map(A1 => n_1691, A2 => n_1703, B1 => new_corner_count(11), B2 => n_1704, Z => n_262);
  g30173 : AO22D0BWP7T port map(A1 => n_1689, A2 => n_1703, B1 => new_corner_count(13), B2 => n_1704, Z => n_261);
  g30174 : AO22D0BWP7T port map(A1 => n_1684, A2 => n_1703, B1 => new_corner_count(18), B2 => n_1704, Z => n_260);
  g30175 : AO22D0BWP7T port map(A1 => n_1683, A2 => n_1703, B1 => new_corner_count(19), B2 => n_1704, Z => n_259);
  g30176 : AO22D0BWP7T port map(A1 => n_1679, A2 => n_1703, B1 => new_corner_count(23), B2 => n_1704, Z => n_258);
  g30177 : AO22D0BWP7T port map(A1 => n_1676, A2 => n_1703, B1 => new_corner_count(26), B2 => n_1704, Z => n_257);
  g30178 : AO22D0BWP7T port map(A1 => n_1675, A2 => n_1703, B1 => new_corner_count(27), B2 => n_1704, Z => n_256);
  g30179 : AO22D0BWP7T port map(A1 => n_1672, A2 => n_1703, B1 => new_corner_count(30), B2 => n_1704, Z => n_255);
  g30180 : NR4D0BWP7T port map(A1 => n_1731, A2 => n_1705, A3 => n_1718, A4 => n_1663, ZN => n_254);
  g30181 : AO22D0BWP7T port map(A1 => n_1685, A2 => n_1703, B1 => new_corner_count(17), B2 => n_1704, Z => n_253);
  g30182 : AO22D0BWP7T port map(A1 => n_1671, A2 => n_1703, B1 => new_corner_count(31), B2 => n_1704, Z => n_252);
  g30183 : MOAI22D0BWP7T port map(A1 => n_151, A2 => n_156, B1 => n_1704, B2 => new_corner_count(1), ZN => n_251);
  g30184 : AO22D0BWP7T port map(A1 => n_1690, A2 => n_1703, B1 => new_corner_count(12), B2 => n_1704, Z => n_250);
  g30185 : AO22D0BWP7T port map(A1 => n_1673, A2 => n_1703, B1 => new_corner_count(29), B2 => n_1704, Z => n_249);
  g30186 : AO22D0BWP7T port map(A1 => n_1681, A2 => n_1703, B1 => new_corner_count(21), B2 => n_1704, Z => n_248);
  g30187 : AO22D0BWP7T port map(A1 => n_1688, A2 => n_1703, B1 => new_corner_count(14), B2 => n_1704, Z => n_247);
  g30188 : AO22D0BWP7T port map(A1 => n_1674, A2 => n_1703, B1 => new_corner_count(28), B2 => n_1704, Z => n_246);
  g30189 : AO22D0BWP7T port map(A1 => n_1677, A2 => n_1703, B1 => new_corner_count(25), B2 => n_1704, Z => n_245);
  g30190 : AO22D0BWP7T port map(A1 => n_1682, A2 => n_1703, B1 => new_corner_count(20), B2 => n_1704, Z => n_244);
  g30191 : AO22D0BWP7T port map(A1 => n_1678, A2 => n_1703, B1 => new_corner_count(24), B2 => n_1704, Z => n_243);
  g30192 : AO22D0BWP7T port map(A1 => n_1687, A2 => n_1703, B1 => new_corner_count(15), B2 => n_1704, Z => n_242);
  g30193 : AO22D0BWP7T port map(A1 => n_1686, A2 => n_1703, B1 => new_corner_count(16), B2 => n_1704, Z => n_241);
  g30194 : NR4D0BWP7T port map(A1 => n_1568, A2 => n_1569, A3 => n_1565, A4 => n_1566, ZN => n_240);
  g30195 : AOI22D0BWP7T port map(A1 => n_152, A2 => n_1179, B1 => N(0), B2 => n_1173, ZN => n_239);
  g30196 : AOI22D0BWP7T port map(A1 => n_153, A2 => n_1161, B1 => N(1), B2 => n_1149, ZN => n_238);
  g30197 : AOI211D0BWP7T port map(A1 => n_1570, A2 => n_1578, B => n_1564, C => n_1567, ZN => n_237);
  g30335 : INVD0BWP7T port map(I => n_228, ZN => n_229);
  g30336 : CKND1BWP7T port map(I => n_225, ZN => n_224);
  g30337 : CKND1BWP7T port map(I => n_217, ZN => n_218);
  g30338 : INVD0BWP7T port map(I => n_214, ZN => n_213);
  g30339 : INVD0BWP7T port map(I => n_212, ZN => n_211);
  g30340 : INVD1BWP7T port map(I => n_208, ZN => n_209);
  g30341 : INVD1BWP7T port map(I => n_206, ZN => n_207);
  g30342 : INVD0BWP7T port map(I => n_205, ZN => n_204);
  g30343 : INVD0BWP7T port map(I => n_203, ZN => n_202);
  g30344 : INVD1BWP7T port map(I => n_195, ZN => n_194);
  g30345 : INVD0BWP7T port map(I => n_193, ZN => n_192);
  g30415 : INR2D0BWP7T port map(A1 => new_N(3), B1 => n_1739, ZN => n_191);
  g30416 : OR2D0BWP7T port map(A1 => n_1739, A2 => new_N(0), Z => n_190);
  g30417 : INR2D0BWP7T port map(A1 => new_N(31), B1 => n_1739, ZN => n_189);
  g30418 : INR2D0BWP7T port map(A1 => new_N(30), B1 => n_1739, ZN => n_188);
  g30419 : NR2D0BWP7T port map(A1 => n_1584, A2 => n_1583, ZN => n_187);
  g30420 : INR2D0BWP7T port map(A1 => new_N(28), B1 => n_1739, ZN => n_186);
  g30421 : INR2D0BWP7T port map(A1 => new_N(27), B1 => n_1739, ZN => n_185);
  g30422 : INR2D0BWP7T port map(A1 => new_N(26), B1 => n_1739, ZN => n_184);
  g30423 : INR2D0BWP7T port map(A1 => new_N(24), B1 => n_1739, ZN => n_183);
  g30424 : INR2D0BWP7T port map(A1 => new_N(29), B1 => n_1739, ZN => n_182);
  g30425 : INR2D0BWP7T port map(A1 => new_N(20), B1 => n_1739, ZN => n_181);
  g30426 : INR2D0BWP7T port map(A1 => new_N(16), B1 => n_1739, ZN => n_180);
  g30427 : INR2D0BWP7T port map(A1 => new_N(19), B1 => n_1739, ZN => n_179);
  g30428 : INR2D0BWP7T port map(A1 => new_N(13), B1 => n_1739, ZN => n_178);
  g30429 : INR2D0BWP7T port map(A1 => new_N(15), B1 => n_1739, ZN => n_177);
  g30430 : INR2D0BWP7T port map(A1 => new_N(18), B1 => n_1739, ZN => n_176);
  g30431 : INR2D0BWP7T port map(A1 => new_N(14), B1 => n_1739, ZN => n_175);
  g30432 : INR2D0BWP7T port map(A1 => new_N(10), B1 => n_1739, ZN => n_174);
  g30433 : INR2D0BWP7T port map(A1 => new_N(7), B1 => n_1739, ZN => n_173);
  g30434 : INR2D0BWP7T port map(A1 => new_N(12), B1 => n_1739, ZN => n_172);
  g30435 : INR2D0BWP7T port map(A1 => new_N(21), B1 => n_1739, ZN => n_171);
  g30436 : INR2D0BWP7T port map(A1 => new_N(6), B1 => n_1739, ZN => n_170);
  g30437 : INR2D0BWP7T port map(A1 => new_N(5), B1 => n_1739, ZN => n_169);
  g30438 : INR2D0BWP7T port map(A1 => new_N(25), B1 => n_1739, ZN => n_168);
  g30439 : INR2D0BWP7T port map(A1 => new_N(11), B1 => n_1739, ZN => n_167);
  g30440 : INR2D0BWP7T port map(A1 => new_N(17), B1 => n_1739, ZN => n_166);
  g30441 : INR2D0BWP7T port map(A1 => new_N(4), B1 => n_1739, ZN => n_165);
  g30442 : ND2D0BWP7T port map(A1 => n_1734, A2 => send_corner_flag, ZN => n_164);
  g30443 : INR2D0BWP7T port map(A1 => new_N(2), B1 => n_1739, ZN => n_163);
  g30444 : INR2D0BWP7T port map(A1 => new_N(1), B1 => n_1739, ZN => n_162);
  g30445 : INR2D0BWP7T port map(A1 => new_N(22), B1 => n_1739, ZN => n_161);
  g30446 : INR2D0BWP7T port map(A1 => new_N(8), B1 => n_1739, ZN => n_160);
  g30447 : INR2D0BWP7T port map(A1 => new_N(9), B1 => n_1739, ZN => n_159);
  g30448 : INR2D0BWP7T port map(A1 => new_N(23), B1 => n_1739, ZN => n_158);
  g30449 : INR2D0BWP7T port map(A1 => n_1654, B1 => n_1650, ZN => n_236);
  g30450 : NR2D0BWP7T port map(A1 => n_1699, A2 => n_1701, ZN => n_235);
  g30451 : NR2D0BWP7T port map(A1 => n_148, A2 => N(3), ZN => n_234);
  g30452 : ND2D0BWP7T port map(A1 => n_1740, A2 => corner_count(1), ZN => n_233);
  g30453 : NR2D0BWP7T port map(A1 => n_1733, A2 => n_1738, ZN => n_232);
  g30454 : NR2D0BWP7T port map(A1 => n_1740, A2 => corner_count(0), ZN => n_231);
  g30455 : ND2D0BWP7T port map(A1 => n_1734, A2 => n_147, ZN => n_230);
  g30456 : NR2D0BWP7T port map(A1 => corner_count(1), A2 => corner_count(2), ZN => n_228);
  g30457 : NR2D0BWP7T port map(A1 => n_1740, A2 => n_146, ZN => n_227);
  g30458 : NR2D0BWP7T port map(A1 => n_148, A2 => N(1), ZN => n_226);
  g30459 : NR2D0BWP7T port map(A1 => n_153, A2 => N(2), ZN => n_225);
  g30460 : NR2D0BWP7T port map(A1 => n_154, A2 => n_149, ZN => n_223);
  g30461 : NR2D0BWP7T port map(A1 => n_1700, A2 => corner_count(0), ZN => n_222);
  g30462 : ND2D0BWP7T port map(A1 => N(2), A2 => N(1), ZN => n_221);
  g30463 : ND2D0BWP7T port map(A1 => n_1700, A2 => n_146, ZN => n_220);
  g30464 : NR2D0BWP7T port map(A1 => N(2), A2 => N(1), ZN => n_219);
  g30465 : ND2D0BWP7T port map(A1 => n_1700, A2 => corner_count(0), ZN => n_217);
  g30466 : ND2D0BWP7T port map(A1 => n_152, A2 => n_153, ZN => n_216);
  g30467 : ND2D0BWP7T port map(A1 => n_148, A2 => n_149, ZN => n_215);
  g30468 : NR2D0BWP7T port map(A1 => n_154, A2 => n_147, ZN => n_214);
  g30469 : NR2D0BWP7T port map(A1 => n_1700, A2 => n_146, ZN => n_212);
  g30470 : ND2D0BWP7T port map(A1 => N(0), A2 => N(1), ZN => n_210);
  g30471 : IND2D0BWP7T port map(A1 => corner_check(5), B1 => n_1653, ZN => n_208);
  g30472 : ND2D0BWP7T port map(A1 => n_1653, A2 => corner_check(5), ZN => n_206);
  g30473 : IND2D0BWP7T port map(A1 => corner_check(5), B1 => n_1732, ZN => n_205);
  g30474 : ND2D0BWP7T port map(A1 => n_1732, A2 => corner_check(5), ZN => n_203);
  g30475 : ND2D0BWP7T port map(A1 => n_1670, A2 => new_tail(1), ZN => n_201);
  g30476 : ND2D0BWP7T port map(A1 => n_1670, A2 => new_tail(2), ZN => n_200);
  g30477 : ND2D0BWP7T port map(A1 => n_1670, A2 => new_tail(0), ZN => n_199);
  g30478 : ND2D0BWP7T port map(A1 => n_1670, A2 => new_tail(3), ZN => n_198);
  g30479 : ND2D0BWP7T port map(A1 => n_1670, A2 => new_tail(5), ZN => n_197);
  g30480 : ND2D0BWP7T port map(A1 => n_1670, A2 => new_tail(4), ZN => n_196);
  g30481 : NR2D0BWP7T port map(A1 => n_1704, A2 => n_1739, ZN => n_195);
  g30482 : NR2D0BWP7T port map(A1 => n_1732, A2 => n_1653, ZN => n_193);
  g30484 : INVD1BWP7T port map(I => reset, ZN => n_157);
  g30485 : INVD0BWP7T port map(I => n_1701, ZN => n_156);
  g30487 : INVD0BWP7T port map(I => n_1734, ZN => n_154);
  g30488 : INVD0BWP7T port map(I => N(1), ZN => n_153);
  g30489 : INVD0BWP7T port map(I => N(0), ZN => n_152);
  g30490 : INVD1BWP7T port map(I => n_1703, ZN => n_151);
  g30492 : CKND1BWP7T port map(I => n_1700, ZN => n_150);
  g30493 : INVD1BWP7T port map(I => N(3), ZN => n_149);
  g30494 : INVD1BWP7T port map(I => N(2), ZN => n_148);
  g30495 : INVD1BWP7T port map(I => N(4), ZN => n_147);
  g30496 : INVD1BWP7T port map(I => corner_count(0), ZN => n_146);
  drc_bufs : INVD4BWP7T port map(I => n_143, ZN => snake_output13(1));
  drc_bufs30498 : INVD1BWP7T port map(I => n_1109, ZN => n_143);
  drc_bufs30500 : INVD4BWP7T port map(I => n_142, ZN => snake_output21(4));
  drc_bufs30502 : INVD1BWP7T port map(I => n_1064, ZN => n_142);
  drc_bufs30504 : INVD4BWP7T port map(I => n_141, ZN => snake_output21(3));
  drc_bufs30506 : INVD1BWP7T port map(I => n_1063, ZN => n_141);
  drc_bufs30508 : INVD4BWP7T port map(I => n_140, ZN => snake_output21(2));
  drc_bufs30510 : INVD1BWP7T port map(I => n_1062, ZN => n_140);
  drc_bufs30512 : INVD4BWP7T port map(I => n_139, ZN => snake_output21(1));
  drc_bufs30514 : INVD1BWP7T port map(I => n_1061, ZN => n_139);
  drc_bufs30516 : INVD4BWP7T port map(I => n_138, ZN => snake_output21(0));
  drc_bufs30518 : INVD1BWP7T port map(I => n_1060, ZN => n_138);
  drc_bufs30520 : INVD4BWP7T port map(I => n_137, ZN => snake_output12(0));
  drc_bufs30522 : INVD1BWP7T port map(I => n_1114, ZN => n_137);
  drc_bufs30524 : INVD4BWP7T port map(I => n_136, ZN => snake_output13(4));
  drc_bufs30526 : INVD1BWP7T port map(I => n_1112, ZN => n_136);
  drc_bufs30528 : INVD4BWP7T port map(I => n_135, ZN => snake_output13(3));
  drc_bufs30530 : INVD1BWP7T port map(I => n_1111, ZN => n_135);
  drc_bufs30532 : INVD4BWP7T port map(I => n_134, ZN => snake_output13(2));
  drc_bufs30534 : INVD1BWP7T port map(I => n_1110, ZN => n_134);
  drc_bufs30536 : INVD4BWP7T port map(I => n_133, ZN => snake_output13(0));
  drc_bufs30538 : INVD1BWP7T port map(I => n_1108, ZN => n_133);
  drc_bufs30540 : INVD4BWP7T port map(I => n_132, ZN => snake_output18(4));
  drc_bufs30542 : INVD1BWP7T port map(I => n_1082, ZN => n_132);
  drc_bufs30544 : INVD4BWP7T port map(I => n_131, ZN => snake_output18(3));
  drc_bufs30546 : INVD1BWP7T port map(I => n_1081, ZN => n_131);
  drc_bufs30548 : INVD4BWP7T port map(I => n_130, ZN => snake_output18(2));
  drc_bufs30550 : INVD1BWP7T port map(I => n_1080, ZN => n_130);
  drc_bufs30552 : INVD4BWP7T port map(I => n_129, ZN => snake_output18(1));
  drc_bufs30554 : INVD1BWP7T port map(I => n_1079, ZN => n_129);
  drc_bufs30556 : INVD4BWP7T port map(I => n_128, ZN => snake_output18(0));
  drc_bufs30558 : INVD1BWP7T port map(I => n_1078, ZN => n_128);
  drc_bufs30560 : INVD4BWP7T port map(I => n_127, ZN => snake_output5(0));
  drc_bufs30562 : INVD1BWP7T port map(I => n_1156, ZN => n_127);
  drc_bufs30564 : INVD4BWP7T port map(I => n_126, ZN => snake_output10(4));
  drc_bufs30566 : INVD1BWP7T port map(I => n_1130, ZN => n_126);
  drc_bufs30568 : INVD4BWP7T port map(I => n_125, ZN => snake_output10(3));
  drc_bufs30570 : INVD1BWP7T port map(I => n_1129, ZN => n_125);
  drc_bufs30572 : INVD4BWP7T port map(I => n_124, ZN => snake_output10(2));
  drc_bufs30574 : INVD1BWP7T port map(I => n_1128, ZN => n_124);
  drc_bufs30576 : INVD4BWP7T port map(I => n_123, ZN => snake_output10(0));
  drc_bufs30578 : INVD1BWP7T port map(I => n_1126, ZN => n_123);
  drc_bufs30580 : INVD4BWP7T port map(I => n_122, ZN => snake_output11(4));
  drc_bufs30582 : INVD1BWP7T port map(I => n_1124, ZN => n_122);
  drc_bufs30584 : INVD4BWP7T port map(I => n_121, ZN => snake_output11(3));
  drc_bufs30586 : INVD1BWP7T port map(I => n_1123, ZN => n_121);
  drc_bufs30588 : INVD4BWP7T port map(I => n_120, ZN => snake_output9(0));
  drc_bufs30590 : INVD1BWP7T port map(I => n_1132, ZN => n_120);
  drc_bufs30592 : INVD4BWP7T port map(I => n_119, ZN => snake_output11(2));
  drc_bufs30594 : INVD1BWP7T port map(I => n_1122, ZN => n_119);
  drc_bufs30596 : INVD4BWP7T port map(I => n_118, ZN => snake_output8(1));
  drc_bufs30598 : INVD1BWP7T port map(I => n_1139, ZN => n_118);
  drc_bufs30600 : INVD4BWP7T port map(I => n_117, ZN => snake_output14(4));
  drc_bufs30602 : INVD1BWP7T port map(I => n_1106, ZN => n_117);
  drc_bufs30604 : INVD4BWP7T port map(I => n_116, ZN => snake_output14(3));
  drc_bufs30606 : INVD1BWP7T port map(I => n_1105, ZN => n_116);
  drc_bufs30608 : INVD4BWP7T port map(I => n_115, ZN => snake_output14(2));
  drc_bufs30610 : INVD1BWP7T port map(I => n_1104, ZN => n_115);
  drc_bufs30612 : INVD4BWP7T port map(I => n_114, ZN => snake_output9(4));
  drc_bufs30614 : INVD1BWP7T port map(I => n_1136, ZN => n_114);
  drc_bufs30616 : INVD4BWP7T port map(I => n_113, ZN => snake_output19(2));
  drc_bufs30618 : INVD1BWP7T port map(I => n_1074, ZN => n_113);
  drc_bufs30620 : INVD4BWP7T port map(I => n_112, ZN => snake_output19(1));
  drc_bufs30622 : INVD1BWP7T port map(I => n_1073, ZN => n_112);
  drc_bufs30624 : INVD4BWP7T port map(I => n_111, ZN => snake_output19(0));
  drc_bufs30626 : INVD1BWP7T port map(I => n_1072, ZN => n_111);
  drc_bufs30628 : INVD4BWP7T port map(I => n_110, ZN => snake_output9(3));
  drc_bufs30630 : INVD1BWP7T port map(I => n_1135, ZN => n_110);
  drc_bufs30632 : INVD4BWP7T port map(I => n_109, ZN => snake_output4(2));
  drc_bufs30634 : INVD1BWP7T port map(I => n_1164, ZN => n_109);
  drc_bufs30636 : INVD4BWP7T port map(I => n_108, ZN => snake_output8(0));
  drc_bufs30638 : INVD1BWP7T port map(I => n_1138, ZN => n_108);
  drc_bufs30640 : INVD4BWP7T port map(I => n_107, ZN => snake_output9(1));
  drc_bufs30642 : INVD1BWP7T port map(I => n_1133, ZN => n_107);
  drc_bufs30644 : INVD4BWP7T port map(I => n_106, ZN => snake_output9(2));
  drc_bufs30646 : INVD1BWP7T port map(I => n_1134, ZN => n_106);
  drc_bufs30648 : INVD4BWP7T port map(I => n_105, ZN => snake_output4(1));
  drc_bufs30650 : INVD1BWP7T port map(I => n_1163, ZN => n_105);
  drc_bufs30652 : INVD4BWP7T port map(I => n_104, ZN => snake_output4(4));
  drc_bufs30654 : INVD1BWP7T port map(I => n_1166, ZN => n_104);
  drc_bufs30656 : INVD4BWP7T port map(I => n_103, ZN => snake_output10(1));
  drc_bufs30658 : INVD1BWP7T port map(I => n_1127, ZN => n_103);
  drc_bufs30660 : INVD4BWP7T port map(I => n_102, ZN => snake_output4(3));
  drc_bufs30662 : INVD1BWP7T port map(I => n_1165, ZN => n_102);
  drc_bufs30664 : INVD4BWP7T port map(I => n_101, ZN => snake_output11(1));
  drc_bufs30666 : INVD1BWP7T port map(I => n_1121, ZN => n_101);
  drc_bufs30668 : INVD4BWP7T port map(I => n_100, ZN => snake_output11(0));
  drc_bufs30670 : INVD1BWP7T port map(I => n_1120, ZN => n_100);
  drc_bufs30672 : INVD4BWP7T port map(I => n_99, ZN => snake_output12(4));
  drc_bufs30674 : INVD1BWP7T port map(I => n_1118, ZN => n_99);
  drc_bufs30676 : INVD4BWP7T port map(I => n_98, ZN => snake_output12(3));
  drc_bufs30678 : INVD1BWP7T port map(I => n_1117, ZN => n_98);
  drc_bufs30680 : INVD4BWP7T port map(I => n_97, ZN => snake_output12(2));
  drc_bufs30682 : INVD1BWP7T port map(I => n_1116, ZN => n_97);
  drc_bufs30684 : INVD4BWP7T port map(I => n_96, ZN => snake_output12(1));
  drc_bufs30686 : INVD1BWP7T port map(I => n_1115, ZN => n_96);
  drc_bufs30688 : INVD4BWP7T port map(I => n_95, ZN => snake_output4(0));
  drc_bufs30690 : INVD1BWP7T port map(I => n_1162, ZN => n_95);
  drc_bufs30692 : INVD4BWP7T port map(I => n_94, ZN => snake_output8(3));
  drc_bufs30694 : INVD1BWP7T port map(I => n_1141, ZN => n_94);
  drc_bufs30696 : INVD4BWP7T port map(I => n_93, ZN => snake_output8(4));
  drc_bufs30698 : INVD1BWP7T port map(I => n_1142, ZN => n_93);
  drc_bufs30700 : INVD4BWP7T port map(I => n_92, ZN => snake_output8(2));
  drc_bufs30702 : INVD1BWP7T port map(I => n_1140, ZN => n_92);
  drc_bufs30704 : INVD4BWP7T port map(I => n_91, ZN => snake_output19(4));
  drc_bufs30706 : INVD1BWP7T port map(I => n_1076, ZN => n_91);
  drc_bufs30708 : INVD4BWP7T port map(I => n_90, ZN => snake_output19(3));
  drc_bufs30710 : INVD1BWP7T port map(I => n_1075, ZN => n_90);
  drc_bufs30712 : INVD4BWP7T port map(I => n_89, ZN => snake_output5(4));
  drc_bufs30714 : INVD1BWP7T port map(I => n_1160, ZN => n_89);
  drc_bufs30716 : INVD4BWP7T port map(I => n_88, ZN => snake_output5(3));
  drc_bufs30718 : INVD1BWP7T port map(I => n_1159, ZN => n_88);
  drc_bufs30720 : INVD4BWP7T port map(I => n_87, ZN => snake_output5(1));
  drc_bufs30722 : INVD1BWP7T port map(I => n_1157, ZN => n_87);
  drc_bufs30724 : INVD4BWP7T port map(I => n_86, ZN => snake_output5(2));
  drc_bufs30726 : INVD1BWP7T port map(I => n_1158, ZN => n_86);
  drc_bufs30728 : INVD4BWP7T port map(I => n_85, ZN => snake_output22(3));
  drc_bufs30730 : INVD1BWP7T port map(I => n_1057, ZN => n_85);
  drc_bufs30732 : INVD4BWP7T port map(I => n_84, ZN => snake_output22(4));
  drc_bufs30734 : INVD1BWP7T port map(I => n_1058, ZN => n_84);
  drc_bufs30736 : INVD4BWP7T port map(I => n_83, ZN => snake_output22(2));
  drc_bufs30738 : INVD1BWP7T port map(I => n_1056, ZN => n_83);
  drc_bufs30740 : INVD4BWP7T port map(I => n_82, ZN => snake_output22(0));
  drc_bufs30742 : INVD1BWP7T port map(I => n_1054, ZN => n_82);
  drc_bufs30744 : INVD4BWP7T port map(I => n_81, ZN => snake_output14(1));
  drc_bufs30746 : INVD1BWP7T port map(I => n_1103, ZN => n_81);
  drc_bufs30748 : INVD4BWP7T port map(I => n_80, ZN => snake_output22(1));
  drc_bufs30750 : INVD1BWP7T port map(I => n_1055, ZN => n_80);
  drc_bufs30752 : INVD4BWP7T port map(I => n_79, ZN => snake_output7(4));
  drc_bufs30754 : INVD1BWP7T port map(I => n_1148, ZN => n_79);
  drc_bufs30756 : INVD4BWP7T port map(I => n_78, ZN => snake_output7(3));
  drc_bufs30758 : INVD1BWP7T port map(I => n_1147, ZN => n_78);
  drc_bufs30760 : INVD4BWP7T port map(I => n_77, ZN => snake_output14(0));
  drc_bufs30762 : INVD1BWP7T port map(I => n_1102, ZN => n_77);
  drc_bufs30764 : INVD4BWP7T port map(I => n_76, ZN => snake_output7(1));
  drc_bufs30766 : INVD1BWP7T port map(I => n_1145, ZN => n_76);
  drc_bufs30768 : INVD4BWP7T port map(I => n_75, ZN => snake_output7(2));
  drc_bufs30770 : INVD1BWP7T port map(I => n_1146, ZN => n_75);
  drc_bufs30772 : INVD4BWP7T port map(I => n_74, ZN => snake_output15(4));
  drc_bufs30774 : INVD1BWP7T port map(I => n_1100, ZN => n_74);
  drc_bufs30776 : INVD4BWP7T port map(I => n_73, ZN => snake_output15(3));
  drc_bufs30778 : INVD1BWP7T port map(I => n_1099, ZN => n_73);
  drc_bufs30780 : INVD4BWP7T port map(I => n_72, ZN => snake_output15(2));
  drc_bufs30782 : INVD1BWP7T port map(I => n_1098, ZN => n_72);
  drc_bufs30784 : INVD4BWP7T port map(I => n_71, ZN => snake_output15(1));
  drc_bufs30786 : INVD1BWP7T port map(I => n_1097, ZN => n_71);
  drc_bufs30788 : INVD4BWP7T port map(I => n_70, ZN => snake_output15(0));
  drc_bufs30790 : INVD1BWP7T port map(I => n_1096, ZN => n_70);
  drc_bufs30792 : INVD4BWP7T port map(I => n_69, ZN => snake_output2(4));
  drc_bufs30794 : INVD1BWP7T port map(I => n_1178, ZN => n_69);
  drc_bufs30796 : INVD4BWP7T port map(I => n_68, ZN => snake_output2(3));
  drc_bufs30798 : INVD1BWP7T port map(I => n_1177, ZN => n_68);
  drc_bufs30800 : INVD4BWP7T port map(I => n_67, ZN => snake_output2(2));
  drc_bufs30802 : INVD1BWP7T port map(I => n_1176, ZN => n_67);
  drc_bufs30804 : INVD4BWP7T port map(I => n_66, ZN => snake_output2(1));
  drc_bufs30806 : INVD1BWP7T port map(I => n_1175, ZN => n_66);
  drc_bufs30808 : INVD4BWP7T port map(I => n_65, ZN => snake_output2(0));
  drc_bufs30810 : INVD1BWP7T port map(I => n_1174, ZN => n_65);
  drc_bufs30812 : INVD4BWP7T port map(I => n_64, ZN => snake_output16(4));
  drc_bufs30814 : INVD1BWP7T port map(I => n_1094, ZN => n_64);
  drc_bufs30816 : INVD4BWP7T port map(I => n_63, ZN => snake_output16(0));
  drc_bufs30818 : INVD1BWP7T port map(I => n_1090, ZN => n_63);
  drc_bufs30820 : INVD4BWP7T port map(I => n_62, ZN => snake_output16(3));
  drc_bufs30822 : INVD1BWP7T port map(I => n_1093, ZN => n_62);
  drc_bufs30824 : INVD4BWP7T port map(I => n_61, ZN => snake_output16(2));
  drc_bufs30826 : INVD1BWP7T port map(I => n_1092, ZN => n_61);
  drc_bufs30828 : INVD4BWP7T port map(I => n_60, ZN => snake_output16(1));
  drc_bufs30830 : INVD1BWP7T port map(I => n_1091, ZN => n_60);
  drc_bufs30832 : INVD4BWP7T port map(I => n_59, ZN => snake_output23(0));
  drc_bufs30834 : INVD1BWP7T port map(I => n_1048, ZN => n_59);
  drc_bufs30836 : INVD4BWP7T port map(I => n_58, ZN => snake_output3(0));
  drc_bufs30838 : INVD1BWP7T port map(I => n_1168, ZN => n_58);
  drc_bufs30840 : INVD4BWP7T port map(I => n_57, ZN => snake_output1(0));
  drc_bufs30842 : INVD1BWP7T port map(I => n_1180, ZN => n_57);
  drc_bufs30844 : INVD4BWP7T port map(I => n_56, ZN => snake_output3(4));
  drc_bufs30846 : INVD1BWP7T port map(I => n_1172, ZN => n_56);
  drc_bufs30848 : INVD4BWP7T port map(I => n_55, ZN => snake_output23(4));
  drc_bufs30850 : INVD1BWP7T port map(I => n_1052, ZN => n_55);
  drc_bufs30852 : INVD4BWP7T port map(I => n_54, ZN => snake_output6(1));
  drc_bufs30854 : INVD1BWP7T port map(I => n_1151, ZN => n_54);
  drc_bufs30856 : INVD4BWP7T port map(I => n_53, ZN => snake_output23(2));
  drc_bufs30858 : INVD1BWP7T port map(I => n_1050, ZN => n_53);
  drc_bufs30860 : INVD4BWP7T port map(I => n_52, ZN => snake_output3(2));
  drc_bufs30862 : INVD1BWP7T port map(I => n_1170, ZN => n_52);
  drc_bufs30864 : INVD4BWP7T port map(I => n_51, ZN => snake_output17(3));
  drc_bufs30866 : INVD1BWP7T port map(I => n_1087, ZN => n_51);
  drc_bufs30868 : INVD4BWP7T port map(I => n_50, ZN => snake_output23(3));
  drc_bufs30870 : INVD1BWP7T port map(I => n_1051, ZN => n_50);
  drc_bufs30872 : INVD4BWP7T port map(I => n_49, ZN => snake_output23(1));
  drc_bufs30874 : INVD1BWP7T port map(I => n_1049, ZN => n_49);
  drc_bufs30876 : INVD4BWP7T port map(I => n_48, ZN => snake_output6(4));
  drc_bufs30878 : INVD1BWP7T port map(I => n_1154, ZN => n_48);
  drc_bufs30880 : INVD4BWP7T port map(I => n_47, ZN => snake_output6(3));
  drc_bufs30882 : INVD1BWP7T port map(I => n_1153, ZN => n_47);
  drc_bufs30884 : INVD4BWP7T port map(I => n_46, ZN => snake_output6(2));
  drc_bufs30886 : INVD1BWP7T port map(I => n_1152, ZN => n_46);
  drc_bufs30888 : INVD4BWP7T port map(I => n_45, ZN => snake_output17(4));
  drc_bufs30890 : INVD1BWP7T port map(I => n_1088, ZN => n_45);
  drc_bufs30892 : INVD4BWP7T port map(I => n_44, ZN => snake_output17(2));
  drc_bufs30894 : INVD1BWP7T port map(I => n_1086, ZN => n_44);
  drc_bufs30896 : INVD4BWP7T port map(I => n_43, ZN => snake_output17(1));
  drc_bufs30898 : INVD1BWP7T port map(I => n_1085, ZN => n_43);
  drc_bufs30900 : INVD4BWP7T port map(I => n_42, ZN => snake_output17(0));
  drc_bufs30902 : INVD1BWP7T port map(I => n_1084, ZN => n_42);
  drc_bufs30904 : INVD4BWP7T port map(I => n_41, ZN => snake_output3(1));
  drc_bufs30906 : INVD1BWP7T port map(I => n_1169, ZN => n_41);
  drc_bufs30908 : INVD4BWP7T port map(I => n_40, ZN => snake_output3(3));
  drc_bufs30910 : INVD1BWP7T port map(I => n_1171, ZN => n_40);
  drc_bufs30912 : INVD4BWP7T port map(I => n_39, ZN => snake_output20(2));
  drc_bufs30914 : INVD1BWP7T port map(I => n_1068, ZN => n_39);
  drc_bufs30916 : INVD4BWP7T port map(I => n_38, ZN => snake_output20(4));
  drc_bufs30918 : INVD1BWP7T port map(I => n_1070, ZN => n_38);
  drc_bufs30920 : INVD4BWP7T port map(I => n_37, ZN => snake_output20(3));
  drc_bufs30922 : INVD1BWP7T port map(I => n_1069, ZN => n_37);
  drc_bufs30924 : INVD4BWP7T port map(I => n_36, ZN => snake_output20(0));
  drc_bufs30926 : INVD1BWP7T port map(I => n_1066, ZN => n_36);
  drc_bufs30928 : INVD4BWP7T port map(I => n_35, ZN => snake_output1(1));
  drc_bufs30930 : INVD1BWP7T port map(I => n_1181, ZN => n_35);
  drc_bufs30932 : INVD4BWP7T port map(I => n_34, ZN => snake_output1(4));
  drc_bufs30934 : INVD1BWP7T port map(I => n_1184, ZN => n_34);
  drc_bufs30936 : INVD4BWP7T port map(I => n_33, ZN => snake_output7(0));
  drc_bufs30938 : INVD1BWP7T port map(I => n_1144, ZN => n_33);
  drc_bufs30940 : INVD4BWP7T port map(I => n_32, ZN => snake_output1(3));
  drc_bufs30942 : INVD1BWP7T port map(I => n_1183, ZN => n_32);
  drc_bufs30944 : INVD4BWP7T port map(I => n_31, ZN => snake_output6(0));
  drc_bufs30946 : INVD1BWP7T port map(I => n_1150, ZN => n_31);
  drc_bufs30948 : INVD4BWP7T port map(I => n_30, ZN => snake_output1(2));
  drc_bufs30950 : INVD1BWP7T port map(I => n_1182, ZN => n_30);
  drc_bufs30952 : INVD4BWP7T port map(I => n_29, ZN => snake_output20(1));
  drc_bufs30954 : INVD1BWP7T port map(I => n_1067, ZN => n_29);
  drc_bufs30956 : INVD4BWP7T port map(I => n_28, ZN => snake_output1(5));
  drc_bufs30958 : INVD1BWP7T port map(I => n_1185, ZN => n_28);
  drc_bufs30961 : INVD4BWP7T port map(I => n_27, ZN => snake_output21(5));
  drc_bufs30962 : INVD1BWP7T port map(I => n_1065, ZN => n_27);
  drc_bufs30965 : INVD4BWP7T port map(I => n_26, ZN => snake_output11(5));
  drc_bufs30966 : INVD1BWP7T port map(I => n_1125, ZN => n_26);
  drc_bufs30969 : INVD4BWP7T port map(I => n_25, ZN => snake_output18(5));
  drc_bufs30970 : INVD1BWP7T port map(I => n_1083, ZN => n_25);
  drc_bufs30973 : INVD4BWP7T port map(I => n_24, ZN => snake_output9(5));
  drc_bufs30974 : INVD1BWP7T port map(I => n_1137, ZN => n_24);
  drc_bufs30977 : INVD4BWP7T port map(I => n_23, ZN => snake_output10(5));
  drc_bufs30978 : INVD1BWP7T port map(I => n_1131, ZN => n_23);
  drc_bufs30981 : INVD4BWP7T port map(I => n_22, ZN => snake_output5(5));
  drc_bufs30982 : INVD1BWP7T port map(I => n_1161, ZN => n_22);
  drc_bufs30985 : INVD4BWP7T port map(I => n_21, ZN => snake_output12(5));
  drc_bufs30986 : INVD1BWP7T port map(I => n_1119, ZN => n_21);
  drc_bufs30989 : INVD4BWP7T port map(I => n_20, ZN => snake_output19(5));
  drc_bufs30990 : INVD1BWP7T port map(I => n_1077, ZN => n_20);
  drc_bufs30993 : INVD4BWP7T port map(I => n_144, ZN => snake_output4(5));
  drc_bufs30994 : INVD1BWP7T port map(I => n_1167, ZN => n_144);
  drc_bufs30997 : INVD4BWP7T port map(I => n_19, ZN => snake_output13(5));
  drc_bufs30998 : INVD1BWP7T port map(I => n_1113, ZN => n_19);
  drc_bufs31001 : INVD4BWP7T port map(I => n_18, ZN => snake_output8(5));
  drc_bufs31002 : INVD1BWP7T port map(I => n_1143, ZN => n_18);
  drc_bufs31005 : INVD4BWP7T port map(I => n_17, ZN => snake_output15(5));
  drc_bufs31006 : INVD1BWP7T port map(I => n_1101, ZN => n_17);
  drc_bufs31009 : INVD4BWP7T port map(I => n_16, ZN => snake_output16(5));
  drc_bufs31010 : INVD1BWP7T port map(I => n_1095, ZN => n_16);
  drc_bufs31013 : INVD4BWP7T port map(I => n_15, ZN => snake_output2(5));
  drc_bufs31014 : INVD1BWP7T port map(I => n_1179, ZN => n_15);
  drc_bufs31017 : INVD4BWP7T port map(I => n_14, ZN => snake_output3(5));
  drc_bufs31018 : INVD1BWP7T port map(I => n_1173, ZN => n_14);
  drc_bufs31021 : INVD4BWP7T port map(I => n_13, ZN => snake_output20(5));
  drc_bufs31022 : INVD1BWP7T port map(I => n_1071, ZN => n_13);
  drc_bufs31025 : INVD4BWP7T port map(I => n_12, ZN => snake_output14(5));
  drc_bufs31026 : INVD1BWP7T port map(I => n_1107, ZN => n_12);
  drc_bufs31029 : INVD4BWP7T port map(I => n_11, ZN => snake_output22(5));
  drc_bufs31030 : INVD1BWP7T port map(I => n_1059, ZN => n_11);
  drc_bufs31033 : INVD4BWP7T port map(I => n_10, ZN => snake_output7(5));
  drc_bufs31034 : INVD1BWP7T port map(I => n_1149, ZN => n_10);
  drc_bufs31037 : INVD4BWP7T port map(I => n_9, ZN => snake_output17(5));
  drc_bufs31038 : INVD1BWP7T port map(I => n_1089, ZN => n_9);
  drc_bufs31041 : INVD4BWP7T port map(I => n_145, ZN => snake_output23(5));
  drc_bufs31042 : INVD1BWP7T port map(I => n_1053, ZN => n_145);
  drc_bufs31045 : INVD4BWP7T port map(I => n_8, ZN => snake_output6(5));
  drc_bufs31046 : INVD1BWP7T port map(I => n_1155, ZN => n_8);
  drc_bufs31049 : INVD4BWP7T port map(I => n_7, ZN => snake_output24(1));
  drc_bufs31050 : INVD1BWP7T port map(I => n_1043, ZN => n_7);
  drc_bufs31053 : INVD4BWP7T port map(I => n_6, ZN => snake_output24(0));
  drc_bufs31054 : INVD1BWP7T port map(I => n_1042, ZN => n_6);
  drc_bufs31057 : INVD4BWP7T port map(I => n_5, ZN => snake_output24(4));
  drc_bufs31058 : INVD1BWP7T port map(I => n_1046, ZN => n_5);
  drc_bufs31061 : INVD4BWP7T port map(I => n_4, ZN => snake_output24(2));
  drc_bufs31062 : INVD1BWP7T port map(I => n_1044, ZN => n_4);
  drc_bufs31065 : INVD4BWP7T port map(I => n_3, ZN => snake_output24(3));
  drc_bufs31066 : INVD1BWP7T port map(I => n_1045, ZN => n_3);
  drc_bufs31069 : INVD4BWP7T port map(I => n_2, ZN => snake_output24(5));
  drc_bufs31070 : INVD1BWP7T port map(I => n_1047, ZN => n_2);
  drc_bufs31072 : BUFFD4BWP7T port map(I => n_1193, Z => snake_list(8));
  drc_bufs31073 : BUFFD4BWP7T port map(I => n_1199, Z => snake_list(14));
  drc_bufs31074 : BUFFD4BWP7T port map(I => n_1188, Z => snake_list(3));
  drc_bufs31075 : BUFFD4BWP7T port map(I => n_1201, Z => snake_list(16));
  drc_bufs31076 : BUFFD4BWP7T port map(I => n_1189, Z => snake_list(4));
  drc_bufs31077 : BUFFD4BWP7T port map(I => n_1187, Z => snake_list(2));
  drc_bufs31078 : BUFFD4BWP7T port map(I => n_1196, Z => snake_list(11));
  drc_bufs31079 : BUFFD4BWP7T port map(I => n_1195, Z => snake_list(10));
  drc_bufs31080 : BUFFD4BWP7T port map(I => n_1186, Z => snake_list(1));
  drc_bufs31081 : BUFFD4BWP7T port map(I => n_1200, Z => snake_list(15));
  drc_bufs31082 : BUFFD4BWP7T port map(I => n_1190, Z => snake_list(5));
  drc_bufs31083 : BUFFD4BWP7T port map(I => n_1198, Z => snake_list(13));
  drc_bufs31084 : BUFFD4BWP7T port map(I => n_1194, Z => snake_list(9));
  drc_bufs31085 : BUFFD4BWP7T port map(I => n_1197, Z => snake_list(12));
  drc_bufs31086 : BUFFD4BWP7T port map(I => n_1191, Z => snake_list(6));
  drc_bufs31087 : BUFFD4BWP7T port map(I => n_1192, Z => snake_list(7));
  g12863 : IND3D1BWP7T port map(A1 => n_610, B1 => n_212, B2 => n_1699, ZN => n_1);
  g31088 : INR3D0BWP7T port map(A1 => n_463, B1 => n_535, B2 => n_429, ZN => n_0);
  g31090 : AO21D0BWP7T port map(A1 => n_1210, A2 => new_corner_flag, B => n_1574, Z => n_1747);
  g31091 : ND3D0BWP7T port map(A1 => n_446, A2 => n_164, A3 => n_240, ZN => n_1748);
  state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => new_state(0), D => n_157, Q => state(0), QN => n_1205);
  state_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => new_state(2), D => n_157, Q => state(2), QN => n_1204);
  g31096 : IND4D0BWP7T port map(A1 => n_1703, B1 => n_1276, B2 => n_1405, B3 => n_1342, ZN => n_1749);
  inc_add_286_38_g321 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_58, A2 => corner_count(31), B1 => inc_add_286_38_n_58, B2 => corner_count(31), ZN => n_1618);
  inc_add_286_38_g322 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_56, A2 => corner_count(30), B1 => inc_add_286_38_n_56, B2 => corner_count(30), ZN => n_1619);
  inc_add_286_38_g323 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_56, B1 => corner_count(30), ZN => inc_add_286_38_n_58);
  inc_add_286_38_g324 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_54, A2 => corner_count(29), B1 => inc_add_286_38_n_54, B2 => corner_count(29), ZN => n_1620);
  inc_add_286_38_g325 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_54, B1 => corner_count(29), ZN => inc_add_286_38_n_56);
  inc_add_286_38_g326 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_52, A2 => corner_count(28), B1 => inc_add_286_38_n_52, B2 => corner_count(28), ZN => n_1621);
  inc_add_286_38_g327 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_52, B1 => corner_count(28), ZN => inc_add_286_38_n_54);
  inc_add_286_38_g328 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_50, A2 => corner_count(27), B1 => inc_add_286_38_n_50, B2 => corner_count(27), ZN => n_1622);
  inc_add_286_38_g329 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_50, B1 => corner_count(27), ZN => inc_add_286_38_n_52);
  inc_add_286_38_g330 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_48, A2 => corner_count(26), B1 => inc_add_286_38_n_48, B2 => corner_count(26), ZN => n_1623);
  inc_add_286_38_g331 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_48, B1 => corner_count(26), ZN => inc_add_286_38_n_50);
  inc_add_286_38_g332 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_46, A2 => corner_count(25), B1 => inc_add_286_38_n_46, B2 => corner_count(25), ZN => n_1624);
  inc_add_286_38_g333 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_46, B1 => corner_count(25), ZN => inc_add_286_38_n_48);
  inc_add_286_38_g334 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_44, A2 => corner_count(24), B1 => inc_add_286_38_n_44, B2 => corner_count(24), ZN => n_1625);
  inc_add_286_38_g335 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_44, B1 => corner_count(24), ZN => inc_add_286_38_n_46);
  inc_add_286_38_g336 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_42, A2 => corner_count(23), B1 => inc_add_286_38_n_42, B2 => corner_count(23), ZN => n_1626);
  inc_add_286_38_g337 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_42, B1 => corner_count(23), ZN => inc_add_286_38_n_44);
  inc_add_286_38_g338 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_40, A2 => corner_count(22), B1 => inc_add_286_38_n_40, B2 => corner_count(22), ZN => n_1627);
  inc_add_286_38_g339 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_40, B1 => corner_count(22), ZN => inc_add_286_38_n_42);
  inc_add_286_38_g340 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_38, A2 => corner_count(21), B1 => inc_add_286_38_n_38, B2 => corner_count(21), ZN => n_1628);
  inc_add_286_38_g341 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_38, B1 => corner_count(21), ZN => inc_add_286_38_n_40);
  inc_add_286_38_g342 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_36, A2 => corner_count(20), B1 => inc_add_286_38_n_36, B2 => corner_count(20), ZN => n_1629);
  inc_add_286_38_g343 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_36, B1 => corner_count(20), ZN => inc_add_286_38_n_38);
  inc_add_286_38_g344 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_34, A2 => corner_count(19), B1 => inc_add_286_38_n_34, B2 => corner_count(19), ZN => n_1630);
  inc_add_286_38_g345 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_34, B1 => corner_count(19), ZN => inc_add_286_38_n_36);
  inc_add_286_38_g346 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_32, A2 => corner_count(18), B1 => inc_add_286_38_n_32, B2 => corner_count(18), ZN => n_1631);
  inc_add_286_38_g347 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_32, B1 => corner_count(18), ZN => inc_add_286_38_n_34);
  inc_add_286_38_g348 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_30, A2 => corner_count(17), B1 => inc_add_286_38_n_30, B2 => corner_count(17), ZN => n_1632);
  inc_add_286_38_g349 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_30, B1 => corner_count(17), ZN => inc_add_286_38_n_32);
  inc_add_286_38_g350 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_28, A2 => corner_count(16), B1 => inc_add_286_38_n_28, B2 => corner_count(16), ZN => n_1633);
  inc_add_286_38_g351 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_28, B1 => corner_count(16), ZN => inc_add_286_38_n_30);
  inc_add_286_38_g352 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_26, A2 => corner_count(15), B1 => inc_add_286_38_n_26, B2 => corner_count(15), ZN => n_1634);
  inc_add_286_38_g353 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_26, B1 => corner_count(15), ZN => inc_add_286_38_n_28);
  inc_add_286_38_g354 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_24, A2 => corner_count(14), B1 => inc_add_286_38_n_24, B2 => corner_count(14), ZN => n_1635);
  inc_add_286_38_g355 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_24, B1 => corner_count(14), ZN => inc_add_286_38_n_26);
  inc_add_286_38_g356 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_22, A2 => corner_count(13), B1 => inc_add_286_38_n_22, B2 => corner_count(13), ZN => n_1636);
  inc_add_286_38_g357 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_22, B1 => corner_count(13), ZN => inc_add_286_38_n_24);
  inc_add_286_38_g358 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_20, A2 => corner_count(12), B1 => inc_add_286_38_n_20, B2 => corner_count(12), ZN => n_1637);
  inc_add_286_38_g359 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_20, B1 => corner_count(12), ZN => inc_add_286_38_n_22);
  inc_add_286_38_g360 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_18, A2 => corner_count(11), B1 => inc_add_286_38_n_18, B2 => corner_count(11), ZN => n_1638);
  inc_add_286_38_g361 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_18, B1 => corner_count(11), ZN => inc_add_286_38_n_20);
  inc_add_286_38_g362 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_16, A2 => corner_count(10), B1 => inc_add_286_38_n_16, B2 => corner_count(10), ZN => n_1639);
  inc_add_286_38_g363 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_16, B1 => corner_count(10), ZN => inc_add_286_38_n_18);
  inc_add_286_38_g364 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_14, A2 => corner_count(9), B1 => inc_add_286_38_n_14, B2 => corner_count(9), ZN => n_1640);
  inc_add_286_38_g365 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_14, B1 => corner_count(9), ZN => inc_add_286_38_n_16);
  inc_add_286_38_g366 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_12, A2 => corner_count(8), B1 => inc_add_286_38_n_12, B2 => corner_count(8), ZN => n_1641);
  inc_add_286_38_g367 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_12, B1 => corner_count(8), ZN => inc_add_286_38_n_14);
  inc_add_286_38_g368 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_10, A2 => corner_count(7), B1 => inc_add_286_38_n_10, B2 => corner_count(7), ZN => n_1642);
  inc_add_286_38_g369 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_10, B1 => corner_count(7), ZN => inc_add_286_38_n_12);
  inc_add_286_38_g370 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_8, A2 => corner_count(6), B1 => inc_add_286_38_n_8, B2 => corner_count(6), ZN => n_1643);
  inc_add_286_38_g371 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_8, B1 => corner_count(6), ZN => inc_add_286_38_n_10);
  inc_add_286_38_g372 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_6, A2 => corner_count(5), B1 => inc_add_286_38_n_6, B2 => corner_count(5), ZN => n_1644);
  inc_add_286_38_g373 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_6, B1 => corner_count(5), ZN => inc_add_286_38_n_8);
  inc_add_286_38_g374 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_4, A2 => corner_count(4), B1 => inc_add_286_38_n_4, B2 => corner_count(4), ZN => n_1645);
  inc_add_286_38_g375 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_4, B1 => corner_count(4), ZN => inc_add_286_38_n_6);
  inc_add_286_38_g376 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_2, A2 => corner_count(3), B1 => inc_add_286_38_n_2, B2 => corner_count(3), ZN => n_1646);
  inc_add_286_38_g377 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_2, B1 => corner_count(3), ZN => inc_add_286_38_n_4);
  inc_add_286_38_g378 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_0, A2 => corner_count(2), B1 => inc_add_286_38_n_0, B2 => corner_count(2), ZN => n_1647);
  inc_add_286_38_g379 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_0, B1 => corner_count(2), ZN => inc_add_286_38_n_2);
  inc_add_286_38_g380 : CKXOR2D0BWP7T port map(A1 => corner_count(0), A2 => corner_count(1), Z => n_1648);
  inc_add_286_38_g381 : ND2D0BWP7T port map(A1 => corner_count(0), A2 => corner_count(1), ZN => inc_add_286_38_n_0);
  inc_add_1070_17_g321 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_58, A2 => N(31), B1 => inc_add_1070_17_n_58, B2 => N(31), ZN => n_1587);
  inc_add_1070_17_g322 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_56, A2 => N(30), B1 => inc_add_1070_17_n_56, B2 => N(30), ZN => n_1588);
  inc_add_1070_17_g323 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_56, B1 => N(30), ZN => inc_add_1070_17_n_58);
  inc_add_1070_17_g324 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_54, A2 => N(29), B1 => inc_add_1070_17_n_54, B2 => N(29), ZN => n_1589);
  inc_add_1070_17_g325 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_54, B1 => N(29), ZN => inc_add_1070_17_n_56);
  inc_add_1070_17_g326 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_52, A2 => N(28), B1 => inc_add_1070_17_n_52, B2 => N(28), ZN => n_1590);
  inc_add_1070_17_g327 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_52, B1 => N(28), ZN => inc_add_1070_17_n_54);
  inc_add_1070_17_g328 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_50, A2 => N(27), B1 => inc_add_1070_17_n_50, B2 => N(27), ZN => n_1591);
  inc_add_1070_17_g329 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_50, B1 => N(27), ZN => inc_add_1070_17_n_52);
  inc_add_1070_17_g330 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_48, A2 => N(26), B1 => inc_add_1070_17_n_48, B2 => N(26), ZN => n_1592);
  inc_add_1070_17_g331 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_48, B1 => N(26), ZN => inc_add_1070_17_n_50);
  inc_add_1070_17_g332 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_46, A2 => N(25), B1 => inc_add_1070_17_n_46, B2 => N(25), ZN => n_1593);
  inc_add_1070_17_g333 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_46, B1 => N(25), ZN => inc_add_1070_17_n_48);
  inc_add_1070_17_g334 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_44, A2 => N(24), B1 => inc_add_1070_17_n_44, B2 => N(24), ZN => n_1594);
  inc_add_1070_17_g335 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_44, B1 => N(24), ZN => inc_add_1070_17_n_46);
  inc_add_1070_17_g336 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_42, A2 => N(23), B1 => inc_add_1070_17_n_42, B2 => N(23), ZN => n_1595);
  inc_add_1070_17_g337 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_42, B1 => N(23), ZN => inc_add_1070_17_n_44);
  inc_add_1070_17_g338 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_40, A2 => N(22), B1 => inc_add_1070_17_n_40, B2 => N(22), ZN => n_1596);
  inc_add_1070_17_g339 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_40, B1 => N(22), ZN => inc_add_1070_17_n_42);
  inc_add_1070_17_g340 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_38, A2 => N(21), B1 => inc_add_1070_17_n_38, B2 => N(21), ZN => n_1597);
  inc_add_1070_17_g341 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_38, B1 => N(21), ZN => inc_add_1070_17_n_40);
  inc_add_1070_17_g342 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_36, A2 => N(20), B1 => inc_add_1070_17_n_36, B2 => N(20), ZN => n_1598);
  inc_add_1070_17_g343 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_36, B1 => N(20), ZN => inc_add_1070_17_n_38);
  inc_add_1070_17_g344 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_34, A2 => N(19), B1 => inc_add_1070_17_n_34, B2 => N(19), ZN => n_1599);
  inc_add_1070_17_g345 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_34, B1 => N(19), ZN => inc_add_1070_17_n_36);
  inc_add_1070_17_g346 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_32, A2 => N(18), B1 => inc_add_1070_17_n_32, B2 => N(18), ZN => n_1600);
  inc_add_1070_17_g347 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_32, B1 => N(18), ZN => inc_add_1070_17_n_34);
  inc_add_1070_17_g348 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_30, A2 => N(17), B1 => inc_add_1070_17_n_30, B2 => N(17), ZN => n_1601);
  inc_add_1070_17_g349 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_30, B1 => N(17), ZN => inc_add_1070_17_n_32);
  inc_add_1070_17_g350 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_28, A2 => N(16), B1 => inc_add_1070_17_n_28, B2 => N(16), ZN => n_1602);
  inc_add_1070_17_g351 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_28, B1 => N(16), ZN => inc_add_1070_17_n_30);
  inc_add_1070_17_g352 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_26, A2 => N(15), B1 => inc_add_1070_17_n_26, B2 => N(15), ZN => n_1603);
  inc_add_1070_17_g353 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_26, B1 => N(15), ZN => inc_add_1070_17_n_28);
  inc_add_1070_17_g354 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_24, A2 => N(14), B1 => inc_add_1070_17_n_24, B2 => N(14), ZN => n_1604);
  inc_add_1070_17_g355 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_24, B1 => N(14), ZN => inc_add_1070_17_n_26);
  inc_add_1070_17_g356 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_22, A2 => N(13), B1 => inc_add_1070_17_n_22, B2 => N(13), ZN => n_1605);
  inc_add_1070_17_g357 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_22, B1 => N(13), ZN => inc_add_1070_17_n_24);
  inc_add_1070_17_g358 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_20, A2 => N(12), B1 => inc_add_1070_17_n_20, B2 => N(12), ZN => n_1606);
  inc_add_1070_17_g359 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_20, B1 => N(12), ZN => inc_add_1070_17_n_22);
  inc_add_1070_17_g360 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_18, A2 => N(11), B1 => inc_add_1070_17_n_18, B2 => N(11), ZN => n_1607);
  inc_add_1070_17_g361 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_18, B1 => N(11), ZN => inc_add_1070_17_n_20);
  inc_add_1070_17_g362 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_16, A2 => N(10), B1 => inc_add_1070_17_n_16, B2 => N(10), ZN => n_1608);
  inc_add_1070_17_g363 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_16, B1 => N(10), ZN => inc_add_1070_17_n_18);
  inc_add_1070_17_g364 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_14, A2 => N(9), B1 => inc_add_1070_17_n_14, B2 => N(9), ZN => n_1609);
  inc_add_1070_17_g365 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_14, B1 => N(9), ZN => inc_add_1070_17_n_16);
  inc_add_1070_17_g366 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_12, A2 => N(8), B1 => inc_add_1070_17_n_12, B2 => N(8), ZN => n_1610);
  inc_add_1070_17_g367 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_12, B1 => N(8), ZN => inc_add_1070_17_n_14);
  inc_add_1070_17_g368 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_10, A2 => N(7), B1 => inc_add_1070_17_n_10, B2 => N(7), ZN => n_1611);
  inc_add_1070_17_g369 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_10, B1 => N(7), ZN => inc_add_1070_17_n_12);
  inc_add_1070_17_g370 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_8, A2 => N(6), B1 => inc_add_1070_17_n_8, B2 => N(6), ZN => n_1612);
  inc_add_1070_17_g371 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_8, B1 => N(6), ZN => inc_add_1070_17_n_10);
  inc_add_1070_17_g372 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_6, A2 => N(5), B1 => inc_add_1070_17_n_6, B2 => N(5), ZN => n_1613);
  inc_add_1070_17_g373 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_6, B1 => N(5), ZN => inc_add_1070_17_n_8);
  inc_add_1070_17_g374 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_4, A2 => N(4), B1 => inc_add_1070_17_n_4, B2 => N(4), ZN => n_1614);
  inc_add_1070_17_g375 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_4, B1 => N(4), ZN => inc_add_1070_17_n_6);
  inc_add_1070_17_g376 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_2, A2 => N(3), B1 => inc_add_1070_17_n_2, B2 => N(3), ZN => n_1615);
  inc_add_1070_17_g377 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_2, B1 => N(3), ZN => inc_add_1070_17_n_4);
  inc_add_1070_17_g378 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_0, A2 => N(2), B1 => inc_add_1070_17_n_0, B2 => N(2), ZN => n_1616);
  inc_add_1070_17_g379 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_0, B1 => N(2), ZN => inc_add_1070_17_n_2);
  inc_add_1070_17_g380 : CKXOR2D0BWP7T port map(A1 => N(0), A2 => N(1), Z => n_1617);
  inc_add_1070_17_g381 : ND2D0BWP7T port map(A1 => N(0), A2 => N(1), ZN => inc_add_1070_17_n_0);
  sub_868_22_g709 : MOAI22D0BWP7T port map(A1 => sub_868_22_n_58, A2 => corner_count(31), B1 => sub_868_22_n_58, B2 => corner_count(31), ZN => n_1671);
  sub_868_22_g710 : IOA21D0BWP7T port map(A1 => sub_868_22_n_56, A2 => corner_count(30), B => sub_868_22_n_58, ZN => n_1672);
  sub_868_22_g711 : OR2D0BWP7T port map(A1 => sub_868_22_n_56, A2 => corner_count(30), Z => sub_868_22_n_58);
  sub_868_22_g712 : IOA21D0BWP7T port map(A1 => sub_868_22_n_54, A2 => corner_count(29), B => sub_868_22_n_56, ZN => n_1673);
  sub_868_22_g713 : OR2D0BWP7T port map(A1 => sub_868_22_n_54, A2 => corner_count(29), Z => sub_868_22_n_56);
  sub_868_22_g714 : IOA21D0BWP7T port map(A1 => sub_868_22_n_52, A2 => corner_count(28), B => sub_868_22_n_54, ZN => n_1674);
  sub_868_22_g715 : OR2D0BWP7T port map(A1 => sub_868_22_n_52, A2 => corner_count(28), Z => sub_868_22_n_54);
  sub_868_22_g716 : IOA21D0BWP7T port map(A1 => sub_868_22_n_50, A2 => corner_count(27), B => sub_868_22_n_52, ZN => n_1675);
  sub_868_22_g717 : OR2D0BWP7T port map(A1 => sub_868_22_n_50, A2 => corner_count(27), Z => sub_868_22_n_52);
  sub_868_22_g718 : IOA21D0BWP7T port map(A1 => sub_868_22_n_48, A2 => corner_count(26), B => sub_868_22_n_50, ZN => n_1676);
  sub_868_22_g719 : OR2D0BWP7T port map(A1 => sub_868_22_n_48, A2 => corner_count(26), Z => sub_868_22_n_50);
  sub_868_22_g720 : IOA21D0BWP7T port map(A1 => sub_868_22_n_46, A2 => corner_count(25), B => sub_868_22_n_48, ZN => n_1677);
  sub_868_22_g721 : OR2D0BWP7T port map(A1 => sub_868_22_n_46, A2 => corner_count(25), Z => sub_868_22_n_48);
  sub_868_22_g722 : IOA21D0BWP7T port map(A1 => sub_868_22_n_44, A2 => corner_count(24), B => sub_868_22_n_46, ZN => n_1678);
  sub_868_22_g723 : OR2D0BWP7T port map(A1 => sub_868_22_n_44, A2 => corner_count(24), Z => sub_868_22_n_46);
  sub_868_22_g724 : IOA21D0BWP7T port map(A1 => sub_868_22_n_42, A2 => corner_count(23), B => sub_868_22_n_44, ZN => n_1679);
  sub_868_22_g725 : OR2D0BWP7T port map(A1 => sub_868_22_n_42, A2 => corner_count(23), Z => sub_868_22_n_44);
  sub_868_22_g726 : IOA21D0BWP7T port map(A1 => sub_868_22_n_40, A2 => corner_count(22), B => sub_868_22_n_42, ZN => n_1680);
  sub_868_22_g727 : OR2D0BWP7T port map(A1 => sub_868_22_n_40, A2 => corner_count(22), Z => sub_868_22_n_42);
  sub_868_22_g728 : IOA21D0BWP7T port map(A1 => sub_868_22_n_38, A2 => corner_count(21), B => sub_868_22_n_40, ZN => n_1681);
  sub_868_22_g729 : OR2D0BWP7T port map(A1 => sub_868_22_n_38, A2 => corner_count(21), Z => sub_868_22_n_40);
  sub_868_22_g730 : IOA21D0BWP7T port map(A1 => sub_868_22_n_36, A2 => corner_count(20), B => sub_868_22_n_38, ZN => n_1682);
  sub_868_22_g731 : OR2D0BWP7T port map(A1 => sub_868_22_n_36, A2 => corner_count(20), Z => sub_868_22_n_38);
  sub_868_22_g732 : IOA21D0BWP7T port map(A1 => sub_868_22_n_34, A2 => corner_count(19), B => sub_868_22_n_36, ZN => n_1683);
  sub_868_22_g733 : OR2D0BWP7T port map(A1 => sub_868_22_n_34, A2 => corner_count(19), Z => sub_868_22_n_36);
  sub_868_22_g734 : IOA21D0BWP7T port map(A1 => sub_868_22_n_32, A2 => corner_count(18), B => sub_868_22_n_34, ZN => n_1684);
  sub_868_22_g735 : OR2D0BWP7T port map(A1 => sub_868_22_n_32, A2 => corner_count(18), Z => sub_868_22_n_34);
  sub_868_22_g736 : IOA21D0BWP7T port map(A1 => sub_868_22_n_30, A2 => corner_count(17), B => sub_868_22_n_32, ZN => n_1685);
  sub_868_22_g737 : OR2D0BWP7T port map(A1 => sub_868_22_n_30, A2 => corner_count(17), Z => sub_868_22_n_32);
  sub_868_22_g738 : IOA21D0BWP7T port map(A1 => sub_868_22_n_28, A2 => corner_count(16), B => sub_868_22_n_30, ZN => n_1686);
  sub_868_22_g739 : OR2D0BWP7T port map(A1 => sub_868_22_n_28, A2 => corner_count(16), Z => sub_868_22_n_30);
  sub_868_22_g740 : IOA21D0BWP7T port map(A1 => sub_868_22_n_26, A2 => corner_count(15), B => sub_868_22_n_28, ZN => n_1687);
  sub_868_22_g741 : OR2D0BWP7T port map(A1 => sub_868_22_n_26, A2 => corner_count(15), Z => sub_868_22_n_28);
  sub_868_22_g742 : IOA21D0BWP7T port map(A1 => sub_868_22_n_24, A2 => corner_count(14), B => sub_868_22_n_26, ZN => n_1688);
  sub_868_22_g743 : OR2D0BWP7T port map(A1 => sub_868_22_n_24, A2 => corner_count(14), Z => sub_868_22_n_26);
  sub_868_22_g744 : IOA21D0BWP7T port map(A1 => sub_868_22_n_22, A2 => corner_count(13), B => sub_868_22_n_24, ZN => n_1689);
  sub_868_22_g745 : OR2D0BWP7T port map(A1 => sub_868_22_n_22, A2 => corner_count(13), Z => sub_868_22_n_24);
  sub_868_22_g746 : IOA21D0BWP7T port map(A1 => sub_868_22_n_20, A2 => corner_count(12), B => sub_868_22_n_22, ZN => n_1690);
  sub_868_22_g747 : OR2D0BWP7T port map(A1 => sub_868_22_n_20, A2 => corner_count(12), Z => sub_868_22_n_22);
  sub_868_22_g748 : IOA21D0BWP7T port map(A1 => sub_868_22_n_18, A2 => corner_count(11), B => sub_868_22_n_20, ZN => n_1691);
  sub_868_22_g749 : OR2D0BWP7T port map(A1 => sub_868_22_n_18, A2 => corner_count(11), Z => sub_868_22_n_20);
  sub_868_22_g750 : IOA21D0BWP7T port map(A1 => sub_868_22_n_16, A2 => corner_count(10), B => sub_868_22_n_18, ZN => n_1692);
  sub_868_22_g751 : OR2D0BWP7T port map(A1 => sub_868_22_n_16, A2 => corner_count(10), Z => sub_868_22_n_18);
  sub_868_22_g752 : IOA21D0BWP7T port map(A1 => sub_868_22_n_14, A2 => corner_count(9), B => sub_868_22_n_16, ZN => n_1693);
  sub_868_22_g753 : OR2D0BWP7T port map(A1 => sub_868_22_n_14, A2 => corner_count(9), Z => sub_868_22_n_16);
  sub_868_22_g754 : IOA21D0BWP7T port map(A1 => sub_868_22_n_12, A2 => corner_count(8), B => sub_868_22_n_14, ZN => n_1694);
  sub_868_22_g755 : OR2D0BWP7T port map(A1 => sub_868_22_n_12, A2 => corner_count(8), Z => sub_868_22_n_14);
  sub_868_22_g756 : IOA21D0BWP7T port map(A1 => sub_868_22_n_10, A2 => corner_count(7), B => sub_868_22_n_12, ZN => n_1695);
  sub_868_22_g757 : OR2D0BWP7T port map(A1 => sub_868_22_n_10, A2 => corner_count(7), Z => sub_868_22_n_12);
  sub_868_22_g758 : IOA21D0BWP7T port map(A1 => sub_868_22_n_8, A2 => corner_count(6), B => sub_868_22_n_10, ZN => n_1696);
  sub_868_22_g759 : OR2D0BWP7T port map(A1 => sub_868_22_n_8, A2 => corner_count(6), Z => sub_868_22_n_10);
  sub_868_22_g760 : IOA21D0BWP7T port map(A1 => sub_868_22_n_6, A2 => corner_count(5), B => sub_868_22_n_8, ZN => n_1697);
  sub_868_22_g761 : OR2D0BWP7T port map(A1 => sub_868_22_n_6, A2 => corner_count(5), Z => sub_868_22_n_8);
  sub_868_22_g762 : IOA21D0BWP7T port map(A1 => sub_868_22_n_4, A2 => corner_count(4), B => sub_868_22_n_6, ZN => n_1698);
  sub_868_22_g763 : OR2D0BWP7T port map(A1 => sub_868_22_n_4, A2 => corner_count(4), Z => sub_868_22_n_6);
  sub_868_22_g764 : IOA21D0BWP7T port map(A1 => sub_868_22_n_2, A2 => corner_count(3), B => sub_868_22_n_4, ZN => n_1699);
  sub_868_22_g765 : OR2D0BWP7T port map(A1 => sub_868_22_n_2, A2 => corner_count(3), Z => sub_868_22_n_4);
  sub_868_22_g766 : IOA21D0BWP7T port map(A1 => sub_868_22_n_0, A2 => corner_count(2), B => sub_868_22_n_2, ZN => n_1700);
  sub_868_22_g767 : OR2D0BWP7T port map(A1 => sub_868_22_n_0, A2 => corner_count(2), Z => sub_868_22_n_2);
  sub_868_22_g768 : IOA21D0BWP7T port map(A1 => corner_count(1), A2 => corner_count(0), B => sub_868_22_n_0, ZN => n_1701);
  sub_868_22_g769 : OR2D0BWP7T port map(A1 => corner_count(0), A2 => corner_count(1), Z => sub_868_22_n_0);
  tie_0_cell : TIELBWP7T port map(ZN => audio(7));

end synthesised;
