configuration or2_behaviour_cfg of or2 is
   for behaviour
   end for;
end or2_behaviour_cfg;
