library IEEE;
use IEEE.std_logic_1164.ALL;

entity rng_tb is
end rng_tb;

