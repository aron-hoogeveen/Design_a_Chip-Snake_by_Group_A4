library IEEE;
use IEEE.std_logic_1164.ALL;

entity itemgenerator_tb is
end itemgenerator_tb;

