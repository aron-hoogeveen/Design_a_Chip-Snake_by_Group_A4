library IEEE;
use IEEE.std_logic_1164.ALL;

entity storage is
   port(clk     				: in  std_logic;
        reset     				: in  std_logic;
	new_head_flag			: in  std_logic;
        new_head  				: in  std_logic_vector(11 downto 0);
	new_corner_flag			: in  std_logic;
        new_corner 				: in  std_logic_vector(5 downto 0);
	new_tail_flag			: in  std_logic;
        new_tail   				: in  std_logic_vector(5 downto 0);
	new_item_set			: in  std_logic;
	remove_item_type			: in  std_logic;
	remove_item_set			: in  std_logic;
	send_corner_flag			: in  std_logic;
        new_item   				: in  std_logic_vector(11 downto 0);
        snake_list 				: out std_logic_vector(16 downto 0);
        item_out_food   				: out std_logic_vector(11 downto 0);
	item_out_power_up			: out std_logic_vector(11 downto 0);
        audio      				: out std_logic_vector(7 downto 0);
	head	   		: out std_logic_vector(11 downto 0);
	tail	   		: out std_logic;
	new_item_clear			: out std_logic;
	clear_head_flag			: out std_logic;
	clear_corner_flag			: out std_logic;
	clear_tail_flag			: out std_logic;
	remove_item_clear			: out std_logic;
	head_send_flag			: out std_logic;
	snake_send_flag			: out std_logic;
	item_send_flag			: out std_logic;
	send_new_corner_clear			: out std_logic;
	snake_output0			: out std_logic_vector(5 downto 0);
	snake_output1			: out std_logic_vector(5 downto 0);
	snake_output2			: out std_logic_vector(5 downto 0);
	snake_output3			: out std_logic_vector(5 downto 0);
	snake_output4			: out std_logic_vector(5 downto 0);
	snake_output5			: out std_logic_vector(5 downto 0);
	snake_output6			: out std_logic_vector(5 downto 0);
	snake_output7			: out std_logic_vector(5 downto 0);
	snake_output8			: out std_logic_vector(5 downto 0);
	snake_output9			: out std_logic_vector(5 downto 0);
	snake_output10			: out std_logic_vector(5 downto 0);
	snake_output11			: out std_logic_vector(5 downto 0);
	snake_output12			: out std_logic_vector(5 downto 0);
	snake_output13			: out std_logic_vector(5 downto 0);
	snake_output14			: out std_logic_vector(5 downto 0);
	snake_output15			: out std_logic_vector(5 downto 0);
	snake_output16			: out std_logic_vector(5 downto 0);
	snake_output17			: out std_logic_vector(5 downto 0);
	snake_output18			: out std_logic_vector(5 downto 0);
	snake_output19			: out std_logic_vector(5 downto 0);
	snake_output20			: out std_logic_vector(5 downto 0);
	snake_output21			: out std_logic_vector(5 downto 0);
	snake_output22			: out std_logic_vector(5 downto 0);
	snake_output23			: out std_logic_vector(5 downto 0);
	snake_output24			: out std_logic_vector(5 downto 0));
	
end storage;

