library IEEE;
use IEEE.std_logic_1164.ALL;

entity v_cnt_control_tb is
end v_cnt_control_tb;

