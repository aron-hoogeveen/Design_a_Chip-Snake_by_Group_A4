library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of and2 is
begin
	z <= a and b;
end behaviour;

