configuration counter4_behaviour_cfg of counter4 is
   for behaviour
   end for;
end counter4_behaviour_cfg;
