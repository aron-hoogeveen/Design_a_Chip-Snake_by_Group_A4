configuration storage_behaviour_storage_cfg of storage is
   for behaviour_storage
   end for;
end storage_behaviour_storage_cfg;
