configuration counter4_routed_cfg of counter4 is
   for routed
   end for;
end counter4_routed_cfg;
