library IEEE;
use IEEE.std_logic_1164.ALL;

entity pulse_speed_tb is
end pulse_speed_tb;

