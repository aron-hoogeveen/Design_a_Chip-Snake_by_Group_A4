library IEEE;
use IEEE.std_logic_1164.ALL;

entity h_counter_tb is
end h_counter_tb;

