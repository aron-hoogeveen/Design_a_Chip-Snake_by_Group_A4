configuration itemgenerator_behaviour_cfg of itemgenerator is
   for behaviour
   end for;
end itemgenerator_behaviour_cfg;
