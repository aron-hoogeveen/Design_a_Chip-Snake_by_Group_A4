library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of xor2 is
begin
	z <= a xor b;
end behaviour;

