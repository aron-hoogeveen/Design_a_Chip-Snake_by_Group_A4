library IEEE;
use IEEE.std_logic_1164.ALL;

entity vga_controller_tb is

end vga_controller_tb;

