library IEEE;
use IEEE.std_logic_1164.ALL;

entity item_image_tb is
end item_image_tb;

