library IEEE;
use IEEE.std_logic_1164.ALL;

entity snake_image_tb is
end snake_image_tb;

