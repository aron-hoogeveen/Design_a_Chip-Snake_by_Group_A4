library IEEE;
use IEEE.std_logic_1164.ALL;

entity color_gen_tb is
end color_gen_tb;

