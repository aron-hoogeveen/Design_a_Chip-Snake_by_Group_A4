library IEEE;
use IEEE.std_logic_1164.ALL;

entity col_detect_tb is
end col_detect_tb;

