configuration rng_routed_cfg of rng is
   for routed
   end for;
end rng_routed_cfg;
