configuration rng_tb_structural_tb of rng_tb is
   for structural
      for all: rng use configuration work.rng_synthesised_cfg;
      end for;
   end for;
end rng_tb_structural_tb;
