configuration counter4_synthesised_cfg of counter4 is
   for synthesised
   end for;
end counter4_synthesised_cfg;
