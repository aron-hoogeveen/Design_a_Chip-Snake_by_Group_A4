library IEEE;
use IEEE.std_logic_1164.ALL;

entity button_react_tb is
end button_react_tb;

