configuration rng_behaviour_cfg of rng is
   for behaviour
   end for;
end rng_behaviour_cfg;
