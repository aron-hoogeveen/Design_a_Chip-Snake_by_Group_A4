library IEEE;
use IEEE.std_logic_1164.ALL;

entity length_tb is
end length_tb;

