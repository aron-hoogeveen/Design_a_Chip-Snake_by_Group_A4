configuration ff_behaviour_cfg of ff is
   for behaviour
   end for;
end ff_behaviour_cfg;
