library IEEE;
use IEEE.std_logic_1164.ALL;

entity inverter is
   port(a : in  std_logic;
        z : out std_logic);
end inverter;

