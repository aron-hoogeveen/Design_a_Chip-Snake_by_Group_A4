library IEEE;
use IEEE.std_logic_1164.ALL;

entity mux is
   port(a : in  std_logic;
        b : in  std_logic;
        x : in  std_logic;
        z : out std_logic);
end mux;

