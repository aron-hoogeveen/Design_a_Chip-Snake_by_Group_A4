library IEEE;
use IEEE.std_logic_1164.ALL;

entity xor2 is
   port(a : in  std_logic;
        b : in  std_logic;
        z : out std_logic);
end xor2;

