library IEEE;
use IEEE.std_logic_1164.ALL;

entity nep_entity is
   port(clk : in  std_logic);
end nep_entity;

