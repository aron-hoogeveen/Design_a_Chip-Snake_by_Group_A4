
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture routed of storage is

  component DEL01BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD6BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD5BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component BUFFD1P5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component CKBD6BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component LHD1BWP7T
    port(D, E : in std_logic; Q, QN : out std_logic);
  end component;

  component LND1BWP7T
    port(D, EN : in std_logic; Q, QN : out std_logic);
  end component;

  component LNQD1BWP7T
    port(D, EN : in std_logic; Q : out std_logic);
  end component;

  component LHQD1BWP7T
    port(D, E : in std_logic; Q : out std_logic);
  end component;

  component IND4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component NR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AO21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component INR4D0BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AN4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component IND3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OR4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; Z : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OA221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IAO21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component OA21D0BWP7T
    port(A1, A2, B : in std_logic; Z : out std_logic);
  end component;

  component ND4D0BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component AOI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component IIND4D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AO22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI211D1BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component CKND1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component OAI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2XD1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component OAI211D0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D2P5BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component NR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component MAOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component CKXOR2D0BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component XNR2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR3D0BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CN, CP, D : in std_logic; Q : out std_logic);
  end component;

  component AO211D0BWP7T
    port(A1, A2, B, C : in std_logic; Z : out std_logic);
  end component;

  component AOI221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; ZN : out std_logic);
  end component;

  component AOI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component IOA21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI222D0BWP7T
    port(A1, A2, B1, B2, C1, C2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI31D0BWP7T
    port(A1, A2, A3, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D1BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AN3D0BWP7T
    port(A1, A2, A3 : in std_logic; Z : out std_logic);
  end component;

  component NR4D1BWP7T
    port(A1, A2, A3, A4 : in std_logic; ZN : out std_logic);
  end component;

  component INR4D1BWP7T
    port(A1, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component AOI33D0BWP7T
    port(A1, A2, A3, B1, B2, B3 : in std_logic; ZN : out std_logic);
  end component;

  component OAI32D0BWP7T
    port(A1, A2, A3, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component HA1D0BWP7T
    port(A, B : in std_logic; CO, S : out std_logic);
  end component;

  component CKND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component IND3D1BWP7T
    port(A1, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CN, CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component TIELBWP7T
    port(ZN : out std_logic);
  end component;

  signal FE_OFN177_n_674, FE_OFN176_n_483, FE_OFN175_snake_list_1, FE_OFN174_snake_list_13, FE_OFN173_snake_list_3 : std_logic;
  signal FE_OFN172_snake_list_10, FE_OFN171_snake_list_5, FE_OFN170_snake_list_15, FE_OFN169_snake_list_8, FE_OFN168_snake_list_2 : std_logic;
  signal FE_OFN167_snake_list_4, FE_OFN166_snake_list_16, FE_OFN165_snake_list_11, FE_OFN164_snake_list_7, FE_OFN163_snake_list_12 : std_logic;
  signal FE_OFN162_snake_list_9, FE_OFN161_snake_list_14, FE_OFN160_snake_list_6, FE_OFN159_snake_output24_5, FE_OFN158_snake_output24_1 : std_logic;
  signal FE_OFN157_snake_output24_2, FE_OFN156_snake_output24_4, FE_OFN155_snake_output24_0, FE_OFN154_snake_output24_3, FE_OFN153_snake_output3_5 : std_logic;
  signal FE_OFN152_snake_output6_5, FE_OFN151_snake_output22_5, FE_OFN150_snake_output7_5, FE_OFN149_snake_output5_5, FE_OFN148_snake_output2_5 : std_logic;
  signal FE_OFN147_snake_output21_5, FE_OFN146_snake_output20_5, FE_OFN145_snake_output15_5, FE_OFN144_snake_output9_5, FE_OFN143_snake_output10_5 : std_logic;
  signal FE_OFN142_snake_output14_5, FE_OFN141_snake_output18_5, FE_OFN140_snake_output12_5, FE_OFN139_snake_output13_5, FE_OFN138_snake_output19_5 : std_logic;
  signal FE_OFN137_snake_output16_5, FE_OFN136_snake_output17_5, FE_OFN135_snake_output11_5, FE_OFN134_snake_output8_5, FE_OFN133_snake_output23_0 : std_logic;
  signal FE_OFN132_snake_output23_3, FE_OFN131_snake_output23_1, FE_OFN130_snake_output23_4, FE_OFN129_snake_output21_3, FE_OFN128_snake_output23_2 : std_logic;
  signal FE_OFN127_snake_output20_3, FE_OFN126_snake_output20_1, FE_OFN125_snake_output22_1, FE_OFN124_snake_output20_0, FE_OFN123_snake_output19_1 : std_logic;
  signal FE_OFN122_snake_output22_3, FE_OFN121_snake_output21_4, FE_OFN120_snake_output21_1, FE_OFN119_snake_output20_4, FE_OFN118_snake_output22_0 : std_logic;
  signal FE_OFN117_snake_output22_4, FE_OFN116_snake_output18_1, FE_OFN115_snake_output18_4, FE_OFN114_snake_output1_2, FE_OFN113_snake_output1_3 : std_logic;
  signal FE_OFN112_snake_output19_3, FE_OFN111_snake_output19_4, FE_OFN110_snake_output20_2, FE_OFN109_snake_output2_2, FE_OFN108_snake_output17_4 : std_logic;
  signal FE_OFN107_snake_output17_3, FE_OFN106_snake_output16_1, FE_OFN105_snake_output5_4, FE_OFN104_snake_output5_3, FE_OFN103_snake_output18_3 : std_logic;
  signal FE_OFN102_snake_output1_1, FE_OFN101_snake_output2_3, FE_OFN100_snake_output21_2, FE_OFN99_snake_output1_0, FE_OFN98_snake_output17_1 : std_logic;
  signal FE_OFN97_snake_output1_4, FE_OFN96_snake_output22_2, FE_OFN95_snake_output7_3, FE_OFN94_snake_output21_0, FE_OFN93_snake_output7_2 : std_logic;
  signal FE_OFN92_snake_output3_2, FE_OFN91_snake_output16_3, FE_OFN90_snake_output19_2, FE_OFN89_snake_output6_0, FE_OFN88_snake_output4_3 : std_logic;
  signal FE_OFN87_snake_output5_2, FE_OFN86_snake_output5_1, FE_OFN85_snake_output2_1, FE_OFN84_snake_output17_0, FE_OFN83_snake_output6_4 : std_logic;
  signal FE_OFN82_snake_output5_0, FE_OFN81_snake_output16_4, FE_OFN80_snake_output3_1, FE_OFN79_snake_output6_3, FE_OFN78_snake_output3_3 : std_logic;
  signal FE_OFN77_snake_output4_2, FE_OFN76_snake_output3_4, FE_OFN75_snake_output4_0, FE_OFN74_snake_output7_0, FE_OFN73_snake_output16_0 : std_logic;
  signal FE_OFN72_snake_output2_0, FE_OFN71_snake_output2_4, FE_OFN70_snake_output7_4, FE_OFN69_snake_output4_4, FE_OFN68_snake_output6_2 : std_logic;
  signal FE_OFN67_snake_output3_0, FE_OFN66_snake_output4_1, FE_OFN65_snake_output12_1, FE_OFN64_snake_output6_1, FE_OFN63_snake_output11_2 : std_logic;
  signal FE_OFN62_snake_output19_0, FE_OFN61_snake_output18_0, FE_OFN60_snake_output12_3, FE_OFN59_snake_output12_2, FE_OFN58_snake_output11_3 : std_logic;
  signal FE_OFN57_snake_output13_2, FE_OFN56_snake_output10_2, FE_OFN55_snake_output11_1, FE_OFN54_snake_output13_3, FE_OFN53_snake_output11_4 : std_logic;
  signal FE_OFN52_snake_output11_0, FE_OFN51_snake_output18_2, FE_OFN50_snake_output15_1, FE_OFN49_snake_output15_2, FE_OFN48_snake_output10_4 : std_logic;
  signal FE_OFN47_snake_output13_1, FE_OFN46_snake_output17_2, FE_OFN45_snake_output9_3, FE_OFN44_snake_output7_1, FE_OFN43_snake_output9_4 : std_logic;
  signal FE_OFN42_snake_output10_0, FE_OFN41_snake_output16_2, FE_OFN40_snake_output12_4, FE_OFN39_snake_output15_3, FE_OFN38_snake_output13_4 : std_logic;
  signal FE_OFN37_snake_output13_0, FE_OFN36_snake_output9_1, FE_OFN35_snake_output9_2, FE_OFN34_snake_output14_1, FE_OFN33_snake_output1_5 : std_logic;
  signal FE_OFN32_snake_output14_2, FE_OFN31_snake_output12_0, FE_OFN30_snake_output10_3, FE_OFN29_snake_output10_1, FE_OFN28_snake_output14_4 : std_logic;
  signal FE_OFN27_snake_output14_0, FE_OFN26_snake_output9_0, FE_OFN25_snake_output8_3, FE_OFN24_snake_output15_4, FE_OFN23_snake_output14_3 : std_logic;
  signal FE_OFN22_snake_output15_0, FE_OFN21_snake_output8_4, FE_OFN20_snake_output8_0, FE_OFN19_snake_output8_1, FE_OFN18_snake_output8_2 : std_logic;
  signal FE_RN_11, FE_OFN6_audio_0, FE_OFN5_audio_0, FE_OFN4_n_1704, FE_OFN3_n_1704 : std_logic;
  signal FE_OFN2_n_1651, FE_OFN1_n_1657, FE_OFN0_n_1657, CTS_6 : std_logic;
  signal new_N : std_logic_vector(31 downto 0);
  signal new_corner_count : std_logic_vector(31 downto 0);
  signal new_state : std_logic_vector(4 downto 0);
  signal corner_count : std_logic_vector(31 downto 0);
  signal N : std_logic_vector(31 downto 0);
  signal state : std_logic_vector(4 downto 0);
  signal corner_check : std_logic_vector(5 downto 0);
  signal shift0 : std_logic_vector(5 downto 0);
  signal shift1 : std_logic_vector(5 downto 0);
  signal shift2 : std_logic_vector(5 downto 0);
  signal shift3 : std_logic_vector(5 downto 0);
  signal shift4 : std_logic_vector(5 downto 0);
  signal shift5 : std_logic_vector(5 downto 0);
  signal shift6 : std_logic_vector(5 downto 0);
  signal shift7 : std_logic_vector(5 downto 0);
  signal shift8 : std_logic_vector(5 downto 0);
  signal shift9 : std_logic_vector(5 downto 0);
  signal shift10 : std_logic_vector(5 downto 0);
  signal shift11 : std_logic_vector(5 downto 0);
  signal shift12 : std_logic_vector(5 downto 0);
  signal shift13 : std_logic_vector(5 downto 0);
  signal shift14 : std_logic_vector(5 downto 0);
  signal shift15 : std_logic_vector(5 downto 0);
  signal shift16 : std_logic_vector(5 downto 0);
  signal shift17 : std_logic_vector(5 downto 0);
  signal shift18 : std_logic_vector(5 downto 0);
  signal shift19 : std_logic_vector(5 downto 0);
  signal shift20 : std_logic_vector(5 downto 0);
  signal shift21 : std_logic_vector(5 downto 0);
  signal shift22 : std_logic_vector(5 downto 0);
  signal shift23 : std_logic_vector(5 downto 0);
  signal UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2, UNCONNECTED3 : std_logic;
  signal UNCONNECTED4, UNCONNECTED5, UNCONNECTED6, UNCONNECTED7, UNCONNECTED8 : std_logic;
  signal UNCONNECTED9, UNCONNECTED10, UNCONNECTED11, UNCONNECTED12, UNCONNECTED13 : std_logic;
  signal UNCONNECTED14, UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18 : std_logic;
  signal UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22, UNCONNECTED23 : std_logic;
  signal UNCONNECTED24, UNCONNECTED25, UNCONNECTED26, UNCONNECTED27, UNCONNECTED28 : std_logic;
  signal UNCONNECTED29, UNCONNECTED30, UNCONNECTED31, UNCONNECTED32, UNCONNECTED33 : std_logic;
  signal UNCONNECTED34, UNCONNECTED35, UNCONNECTED36, UNCONNECTED37, UNCONNECTED38 : std_logic;
  signal UNCONNECTED39, UNCONNECTED40, UNCONNECTED41, UNCONNECTED42, inc_add_286_38_n_0 : std_logic;
  signal inc_add_286_38_n_2, inc_add_286_38_n_4, inc_add_286_38_n_6, inc_add_286_38_n_8, inc_add_286_38_n_10 : std_logic;
  signal inc_add_286_38_n_12, inc_add_286_38_n_14, inc_add_286_38_n_16, inc_add_286_38_n_18, inc_add_286_38_n_20 : std_logic;
  signal inc_add_286_38_n_22, inc_add_286_38_n_24, inc_add_286_38_n_26, inc_add_286_38_n_28, inc_add_286_38_n_30 : std_logic;
  signal inc_add_286_38_n_32, inc_add_286_38_n_34, inc_add_286_38_n_36, inc_add_286_38_n_38, inc_add_286_38_n_40 : std_logic;
  signal inc_add_286_38_n_42, inc_add_286_38_n_44, inc_add_286_38_n_46, inc_add_286_38_n_48, inc_add_286_38_n_50 : std_logic;
  signal inc_add_286_38_n_52, inc_add_286_38_n_54, inc_add_286_38_n_56, inc_add_286_38_n_58, inc_add_1070_17_n_0 : std_logic;
  signal inc_add_1070_17_n_2, inc_add_1070_17_n_4, inc_add_1070_17_n_6, inc_add_1070_17_n_8, inc_add_1070_17_n_10 : std_logic;
  signal inc_add_1070_17_n_12, inc_add_1070_17_n_14, inc_add_1070_17_n_16, inc_add_1070_17_n_18, inc_add_1070_17_n_20 : std_logic;
  signal inc_add_1070_17_n_22, inc_add_1070_17_n_24, inc_add_1070_17_n_26, inc_add_1070_17_n_28, inc_add_1070_17_n_30 : std_logic;
  signal inc_add_1070_17_n_32, inc_add_1070_17_n_34, inc_add_1070_17_n_36, inc_add_1070_17_n_38, inc_add_1070_17_n_40 : std_logic;
  signal inc_add_1070_17_n_42, inc_add_1070_17_n_44, inc_add_1070_17_n_46, inc_add_1070_17_n_48, inc_add_1070_17_n_50 : std_logic;
  signal inc_add_1070_17_n_52, inc_add_1070_17_n_54, inc_add_1070_17_n_56, inc_add_1070_17_n_58, n_0 : std_logic;
  signal n_1, n_144, n_145, n_146, n_147 : std_logic;
  signal n_148, n_149, n_150, n_151, n_152 : std_logic;
  signal n_153, n_154, n_155, n_156, n_157 : std_logic;
  signal n_158, n_159, n_160, n_161, n_162 : std_logic;
  signal n_163, n_164, n_165, n_166, n_167 : std_logic;
  signal n_168, n_169, n_170, n_171, n_172 : std_logic;
  signal n_173, n_174, n_175, n_176, n_177 : std_logic;
  signal n_178, n_179, n_180, n_181, n_182 : std_logic;
  signal n_183, n_184, n_185, n_186, n_187 : std_logic;
  signal n_188, n_189, n_190, n_191, n_192 : std_logic;
  signal n_193, n_194, n_195, n_196, n_197 : std_logic;
  signal n_198, n_199, n_200, n_201, n_202 : std_logic;
  signal n_203, n_204, n_205, n_206, n_207 : std_logic;
  signal n_208, n_209, n_210, n_211, n_212 : std_logic;
  signal n_213, n_214, n_215, n_216, n_217 : std_logic;
  signal n_218, n_219, n_220, n_221, n_222 : std_logic;
  signal n_223, n_224, n_225, n_226, n_227 : std_logic;
  signal n_228, n_229, n_230, n_231, n_232 : std_logic;
  signal n_233, n_234, n_235, n_236, n_237 : std_logic;
  signal n_238, n_239, n_240, n_241, n_242 : std_logic;
  signal n_243, n_244, n_245, n_246, n_247 : std_logic;
  signal n_248, n_249, n_250, n_251, n_252 : std_logic;
  signal n_253, n_254, n_255, n_256, n_257 : std_logic;
  signal n_258, n_259, n_260, n_261, n_262 : std_logic;
  signal n_263, n_264, n_265, n_266, n_267 : std_logic;
  signal n_268, n_269, n_270, n_271, n_272 : std_logic;
  signal n_273, n_274, n_275, n_276, n_277 : std_logic;
  signal n_278, n_279, n_280, n_281, n_282 : std_logic;
  signal n_283, n_284, n_285, n_286, n_287 : std_logic;
  signal n_288, n_289, n_290, n_291, n_292 : std_logic;
  signal n_293, n_294, n_295, n_296, n_297 : std_logic;
  signal n_298, n_299, n_300, n_301, n_302 : std_logic;
  signal n_303, n_304, n_305, n_306, n_307 : std_logic;
  signal n_308, n_309, n_310, n_311, n_312 : std_logic;
  signal n_313, n_314, n_315, n_316, n_317 : std_logic;
  signal n_318, n_319, n_320, n_321, n_322 : std_logic;
  signal n_323, n_324, n_325, n_326, n_327 : std_logic;
  signal n_328, n_329, n_330, n_331, n_332 : std_logic;
  signal n_333, n_334, n_335, n_336, n_337 : std_logic;
  signal n_338, n_339, n_340, n_341, n_342 : std_logic;
  signal n_343, n_344, n_345, n_346, n_347 : std_logic;
  signal n_348, n_349, n_350, n_351, n_352 : std_logic;
  signal n_353, n_354, n_355, n_356, n_357 : std_logic;
  signal n_358, n_359, n_360, n_361, n_362 : std_logic;
  signal n_363, n_364, n_365, n_366, n_367 : std_logic;
  signal n_368, n_369, n_370, n_371, n_372 : std_logic;
  signal n_373, n_374, n_375, n_376, n_377 : std_logic;
  signal n_378, n_379, n_380, n_381, n_382 : std_logic;
  signal n_383, n_384, n_385, n_386, n_387 : std_logic;
  signal n_388, n_389, n_390, n_391, n_392 : std_logic;
  signal n_393, n_394, n_395, n_396, n_397 : std_logic;
  signal n_398, n_399, n_400, n_401, n_402 : std_logic;
  signal n_403, n_404, n_405, n_406, n_407 : std_logic;
  signal n_408, n_409, n_410, n_411, n_412 : std_logic;
  signal n_413, n_414, n_415, n_416, n_417 : std_logic;
  signal n_418, n_419, n_420, n_421, n_422 : std_logic;
  signal n_423, n_424, n_425, n_426, n_427 : std_logic;
  signal n_428, n_429, n_430, n_431, n_432 : std_logic;
  signal n_433, n_434, n_435, n_436, n_437 : std_logic;
  signal n_438, n_439, n_440, n_441, n_442 : std_logic;
  signal n_443, n_444, n_445, n_446, n_447 : std_logic;
  signal n_448, n_449, n_450, n_451, n_452 : std_logic;
  signal n_453, n_454, n_455, n_456, n_457 : std_logic;
  signal n_458, n_459, n_460, n_461, n_462 : std_logic;
  signal n_463, n_464, n_465, n_466, n_467 : std_logic;
  signal n_468, n_469, n_470, n_471, n_472 : std_logic;
  signal n_473, n_474, n_475, n_476, n_477 : std_logic;
  signal n_478, n_479, n_480, n_481, n_482 : std_logic;
  signal n_483, n_484, n_485, n_486, n_487 : std_logic;
  signal n_488, n_489, n_490, n_491, n_492 : std_logic;
  signal n_493, n_494, n_495, n_496, n_497 : std_logic;
  signal n_498, n_499, n_500, n_501, n_502 : std_logic;
  signal n_503, n_504, n_505, n_506, n_507 : std_logic;
  signal n_508, n_509, n_510, n_511, n_512 : std_logic;
  signal n_513, n_514, n_515, n_516, n_517 : std_logic;
  signal n_518, n_519, n_520, n_521, n_522 : std_logic;
  signal n_523, n_524, n_525, n_526, n_527 : std_logic;
  signal n_528, n_529, n_530, n_531, n_532 : std_logic;
  signal n_533, n_534, n_535, n_536, n_537 : std_logic;
  signal n_538, n_539, n_540, n_541, n_542 : std_logic;
  signal n_543, n_544, n_545, n_546, n_547 : std_logic;
  signal n_549, n_550, n_551, n_552, n_553 : std_logic;
  signal n_554, n_555, n_556, n_557, n_558 : std_logic;
  signal n_559, n_560, n_561, n_562, n_563 : std_logic;
  signal n_564, n_565, n_566, n_567, n_568 : std_logic;
  signal n_569, n_570, n_571, n_572, n_573 : std_logic;
  signal n_574, n_575, n_576, n_577, n_578 : std_logic;
  signal n_579, n_580, n_581, n_582, n_583 : std_logic;
  signal n_584, n_585, n_586, n_587, n_588 : std_logic;
  signal n_589, n_590, n_591, n_592, n_593 : std_logic;
  signal n_594, n_595, n_596, n_597, n_598 : std_logic;
  signal n_599, n_600, n_601, n_602, n_603 : std_logic;
  signal n_604, n_605, n_606, n_607, n_608 : std_logic;
  signal n_609, n_610, n_611, n_612, n_613 : std_logic;
  signal n_614, n_615, n_616, n_617, n_618 : std_logic;
  signal n_619, n_620, n_621, n_622, n_623 : std_logic;
  signal n_624, n_625, n_626, n_627, n_628 : std_logic;
  signal n_629, n_630, n_631, n_632, n_633 : std_logic;
  signal n_634, n_635, n_636, n_637, n_638 : std_logic;
  signal n_639, n_640, n_641, n_642, n_643 : std_logic;
  signal n_644, n_645, n_646, n_647, n_648 : std_logic;
  signal n_649, n_650, n_651, n_652, n_653 : std_logic;
  signal n_654, n_655, n_656, n_657, n_658 : std_logic;
  signal n_659, n_660, n_661, n_662, n_663 : std_logic;
  signal n_664, n_665, n_666, n_667, n_668 : std_logic;
  signal n_669, n_670, n_671, n_672, n_673 : std_logic;
  signal n_674, n_675, n_676, n_677, n_678 : std_logic;
  signal n_679, n_680, n_681, n_682, n_683 : std_logic;
  signal n_684, n_685, n_686, n_687, n_688 : std_logic;
  signal n_689, n_690, n_691, n_692, n_693 : std_logic;
  signal n_694, n_695, n_696, n_697, n_698 : std_logic;
  signal n_699, n_700, n_701, n_702, n_703 : std_logic;
  signal n_704, n_705, n_706, n_707, n_708 : std_logic;
  signal n_709, n_710, n_711, n_712, n_713 : std_logic;
  signal n_714, n_715, n_716, n_717, n_718 : std_logic;
  signal n_719, n_720, n_721, n_722, n_723 : std_logic;
  signal n_724, n_725, n_726, n_727, n_728 : std_logic;
  signal n_729, n_730, n_731, n_732, n_733 : std_logic;
  signal n_734, n_735, n_736, n_737, n_738 : std_logic;
  signal n_739, n_740, n_741, n_742, n_743 : std_logic;
  signal n_744, n_745, n_746, n_747, n_748 : std_logic;
  signal n_749, n_750, n_751, n_752, n_753 : std_logic;
  signal n_754, n_755, n_756, n_757, n_758 : std_logic;
  signal n_759, n_760, n_761, n_762, n_763 : std_logic;
  signal n_764, n_765, n_766, n_767, n_768 : std_logic;
  signal n_769, n_770, n_771, n_772, n_773 : std_logic;
  signal n_774, n_775, n_776, n_777, n_778 : std_logic;
  signal n_779, n_780, n_781, n_782, n_783 : std_logic;
  signal n_784, n_785, n_786, n_787, n_788 : std_logic;
  signal n_789, n_790, n_791, n_792, n_793 : std_logic;
  signal n_794, n_795, n_796, n_797, n_798 : std_logic;
  signal n_799, n_800, n_801, n_802, n_803 : std_logic;
  signal n_804, n_805, n_806, n_807, n_808 : std_logic;
  signal n_809, n_810, n_811, n_812, n_813 : std_logic;
  signal n_814, n_815, n_816, n_817, n_818 : std_logic;
  signal n_819, n_820, n_821, n_822, n_823 : std_logic;
  signal n_824, n_825, n_826, n_827, n_828 : std_logic;
  signal n_829, n_830, n_831, n_832, n_833 : std_logic;
  signal n_834, n_835, n_836, n_837, n_838 : std_logic;
  signal n_839, n_840, n_841, n_842, n_843 : std_logic;
  signal n_844, n_845, n_846, n_847, n_848 : std_logic;
  signal n_849, n_850, n_851, n_852, n_853 : std_logic;
  signal n_854, n_855, n_856, n_857, n_858 : std_logic;
  signal n_859, n_860, n_861, n_862, n_863 : std_logic;
  signal n_864, n_865, n_866, n_867, n_868 : std_logic;
  signal n_869, n_870, n_871, n_872, n_873 : std_logic;
  signal n_874, n_875, n_876, n_877, n_878 : std_logic;
  signal n_879, n_880, n_881, n_882, n_883 : std_logic;
  signal n_884, n_885, n_886, n_887, n_888 : std_logic;
  signal n_889, n_890, n_891, n_892, n_893 : std_logic;
  signal n_894, n_895, n_896, n_897, n_898 : std_logic;
  signal n_899, n_900, n_901, n_902, n_903 : std_logic;
  signal n_904, n_905, n_906, n_907, n_908 : std_logic;
  signal n_909, n_910, n_911, n_912, n_913 : std_logic;
  signal n_914, n_915, n_916, n_917, n_918 : std_logic;
  signal n_919, n_920, n_921, n_922, n_923 : std_logic;
  signal n_924, n_925, n_926, n_927, n_928 : std_logic;
  signal n_929, n_930, n_931, n_932, n_933 : std_logic;
  signal n_934, n_935, n_936, n_937, n_938 : std_logic;
  signal n_939, n_940, n_941, n_942, n_943 : std_logic;
  signal n_944, n_945, n_946, n_947, n_948 : std_logic;
  signal n_949, n_950, n_951, n_952, n_953 : std_logic;
  signal n_954, n_955, n_956, n_957, n_958 : std_logic;
  signal n_959, n_960, n_961, n_962, n_963 : std_logic;
  signal n_964, n_965, n_966, n_967, n_968 : std_logic;
  signal n_969, n_970, n_971, n_972, n_973 : std_logic;
  signal n_974, n_975, n_976, n_977, n_978 : std_logic;
  signal n_979, n_980, n_981, n_982, n_983 : std_logic;
  signal n_984, n_985, n_986, n_987, n_988 : std_logic;
  signal n_989, n_990, n_991, n_992, n_993 : std_logic;
  signal n_994, n_995, n_996, n_997, n_998 : std_logic;
  signal n_999, n_1000, n_1001, n_1002, n_1003 : std_logic;
  signal n_1004, n_1005, n_1006, n_1007, n_1008 : std_logic;
  signal n_1009, n_1010, n_1011, n_1012, n_1013 : std_logic;
  signal n_1014, n_1015, n_1016, n_1017, n_1018 : std_logic;
  signal n_1019, n_1020, n_1021, n_1022, n_1023 : std_logic;
  signal n_1024, n_1025, n_1026, n_1027, n_1028 : std_logic;
  signal n_1029, n_1030, n_1031, n_1032, n_1033 : std_logic;
  signal n_1034, n_1035, n_1036, n_1037, n_1038 : std_logic;
  signal n_1039, n_1040, n_1041, n_1053, n_1167 : std_logic;
  signal n_1202, n_1203, n_1204, n_1205, n_1206 : std_logic;
  signal n_1207, n_1208, n_1209, n_1210, n_1211 : std_logic;
  signal n_1212, n_1214, n_1215, n_1216, n_1217 : std_logic;
  signal n_1218, n_1219, n_1220, n_1221, n_1222 : std_logic;
  signal n_1223, n_1224, n_1225, n_1226, n_1227 : std_logic;
  signal n_1228, n_1229, n_1230, n_1231, n_1232 : std_logic;
  signal n_1233, n_1234, n_1235, n_1236, n_1237 : std_logic;
  signal n_1238, n_1239, n_1240, n_1241, n_1242 : std_logic;
  signal n_1243, n_1244, n_1245, n_1246, n_1247 : std_logic;
  signal n_1248, n_1249, n_1250, n_1251, n_1252 : std_logic;
  signal n_1253, n_1254, n_1255, n_1256, n_1257 : std_logic;
  signal n_1258, n_1259, n_1260, n_1261, n_1262 : std_logic;
  signal n_1263, n_1264, n_1265, n_1266, n_1267 : std_logic;
  signal n_1268, n_1269, n_1270, n_1271, n_1272 : std_logic;
  signal n_1273, n_1274, n_1275, n_1276, n_1277 : std_logic;
  signal n_1278, n_1279, n_1280, n_1281, n_1282 : std_logic;
  signal n_1283, n_1284, n_1285, n_1286, n_1287 : std_logic;
  signal n_1288, n_1289, n_1290, n_1291, n_1292 : std_logic;
  signal n_1293, n_1294, n_1295, n_1296, n_1297 : std_logic;
  signal n_1298, n_1299, n_1300, n_1301, n_1302 : std_logic;
  signal n_1303, n_1304, n_1305, n_1306, n_1307 : std_logic;
  signal n_1309, n_1310, n_1311, n_1312, n_1313 : std_logic;
  signal n_1314, n_1315, n_1316, n_1317, n_1318 : std_logic;
  signal n_1319, n_1320, n_1321, n_1322, n_1323 : std_logic;
  signal n_1324, n_1325, n_1326, n_1327, n_1328 : std_logic;
  signal n_1329, n_1330, n_1331, n_1332, n_1333 : std_logic;
  signal n_1334, n_1335, n_1336, n_1337, n_1338 : std_logic;
  signal n_1339, n_1340, n_1341, n_1342, n_1343 : std_logic;
  signal n_1344, n_1345, n_1346, n_1347, n_1348 : std_logic;
  signal n_1349, n_1350, n_1351, n_1352, n_1353 : std_logic;
  signal n_1354, n_1355, n_1357, n_1358, n_1359 : std_logic;
  signal n_1360, n_1361, n_1362, n_1363, n_1364 : std_logic;
  signal n_1365, n_1366, n_1367, n_1368, n_1369 : std_logic;
  signal n_1370, n_1371, n_1372, n_1373, n_1374 : std_logic;
  signal n_1375, n_1376, n_1377, n_1378, n_1379 : std_logic;
  signal n_1380, n_1381, n_1382, n_1383, n_1384 : std_logic;
  signal n_1385, n_1386, n_1387, n_1388, n_1389 : std_logic;
  signal n_1390, n_1391, n_1392, n_1393, n_1394 : std_logic;
  signal n_1395, n_1396, n_1397, n_1399, n_1400 : std_logic;
  signal n_1401, n_1402, n_1403, n_1404, n_1405 : std_logic;
  signal n_1406, n_1407, n_1408, n_1409, n_1410 : std_logic;
  signal n_1411, n_1413, n_1414, n_1415, n_1416 : std_logic;
  signal n_1417, n_1418, n_1419, n_1420, n_1421 : std_logic;
  signal n_1422, n_1423, n_1424, n_1425, n_1426 : std_logic;
  signal n_1564, n_1565, n_1566, n_1567, n_1568 : std_logic;
  signal n_1569, n_1570, n_1571, n_1572, n_1573 : std_logic;
  signal n_1574, n_1575, n_1578, n_1579, n_1580 : std_logic;
  signal n_1581, n_1582, n_1583, n_1584, n_1585 : std_logic;
  signal n_1587, n_1588, n_1589, n_1590, n_1591 : std_logic;
  signal n_1592, n_1593, n_1594, n_1595, n_1596 : std_logic;
  signal n_1597, n_1598, n_1599, n_1600, n_1601 : std_logic;
  signal n_1602, n_1603, n_1604, n_1605, n_1606 : std_logic;
  signal n_1607, n_1608, n_1609, n_1610, n_1611 : std_logic;
  signal n_1612, n_1613, n_1614, n_1615, n_1616 : std_logic;
  signal n_1617, n_1618, n_1619, n_1620, n_1621 : std_logic;
  signal n_1622, n_1623, n_1624, n_1625, n_1626 : std_logic;
  signal n_1627, n_1628, n_1629, n_1630, n_1631 : std_logic;
  signal n_1632, n_1633, n_1634, n_1635, n_1636 : std_logic;
  signal n_1637, n_1638, n_1639, n_1640, n_1641 : std_logic;
  signal n_1642, n_1643, n_1644, n_1645, n_1646 : std_logic;
  signal n_1647, n_1648, n_1649, n_1650, n_1651 : std_logic;
  signal n_1652, n_1653, n_1654, n_1657, n_1662 : std_logic;
  signal n_1663, n_1670, n_1671, n_1672, n_1673 : std_logic;
  signal n_1674, n_1675, n_1676, n_1677, n_1678 : std_logic;
  signal n_1679, n_1680, n_1681, n_1682, n_1683 : std_logic;
  signal n_1684, n_1685, n_1686, n_1687, n_1688 : std_logic;
  signal n_1689, n_1690, n_1691, n_1692, n_1693 : std_logic;
  signal n_1694, n_1695, n_1696, n_1697, n_1698 : std_logic;
  signal n_1699, n_1700, n_1701, n_1703, n_1704 : std_logic;
  signal n_1705, n_1718, n_1731, n_1732, n_1733 : std_logic;
  signal n_1734, n_1735, n_1736, n_1737, n_1738 : std_logic;
  signal n_1739, n_1740, n_1742, n_1747, n_1748 : std_logic;
  signal n_1749, sub_868_22_n_0, sub_868_22_n_2, sub_868_22_n_4, sub_868_22_n_6 : std_logic;
  signal sub_868_22_n_8, sub_868_22_n_10, sub_868_22_n_12, sub_868_22_n_14, sub_868_22_n_16 : std_logic;
  signal sub_868_22_n_18, sub_868_22_n_20, sub_868_22_n_22, sub_868_22_n_24, sub_868_22_n_26 : std_logic;
  signal sub_868_22_n_28, sub_868_22_n_30, sub_868_22_n_32, sub_868_22_n_34, sub_868_22_n_36 : std_logic;
  signal sub_868_22_n_38, sub_868_22_n_40, sub_868_22_n_42, sub_868_22_n_44, sub_868_22_n_46 : std_logic;
  signal sub_868_22_n_48, sub_868_22_n_50, sub_868_22_n_52, sub_868_22_n_54, sub_868_22_n_56 : std_logic;
  signal sub_868_22_n_58 : std_logic;

begin

  audio(0) <= FE_RN_11;
  FE_OFC177_n_674 : DEL01BWP7T port map(I => n_674, Z => FE_OFN177_n_674);
  FE_OFC176_n_483 : DEL01BWP7T port map(I => n_483, Z => FE_OFN176_n_483);
  FE_OFC175_snake_list_1 : BUFFD5BWP7T port map(I => FE_OFN175_snake_list_1, Z => snake_list(1));
  FE_OFC174_snake_list_13 : BUFFD5BWP7T port map(I => FE_OFN174_snake_list_13, Z => snake_list(13));
  FE_OFC173_snake_list_3 : BUFFD5BWP7T port map(I => FE_OFN173_snake_list_3, Z => snake_list(3));
  FE_OFC172_snake_list_10 : BUFFD5BWP7T port map(I => FE_OFN172_snake_list_10, Z => snake_list(10));
  FE_OFC171_snake_list_5 : BUFFD5BWP7T port map(I => FE_OFN171_snake_list_5, Z => snake_list(5));
  FE_OFC170_snake_list_15 : BUFFD5BWP7T port map(I => FE_OFN170_snake_list_15, Z => snake_list(15));
  FE_OFC169_snake_list_8 : BUFFD5BWP7T port map(I => FE_OFN169_snake_list_8, Z => snake_list(8));
  FE_OFC168_snake_list_2 : BUFFD5BWP7T port map(I => FE_OFN168_snake_list_2, Z => snake_list(2));
  FE_OFC167_snake_list_4 : BUFFD5BWP7T port map(I => FE_OFN167_snake_list_4, Z => snake_list(4));
  FE_OFC166_snake_list_16 : BUFFD5BWP7T port map(I => FE_OFN166_snake_list_16, Z => snake_list(16));
  FE_OFC165_snake_list_11 : BUFFD5BWP7T port map(I => FE_OFN165_snake_list_11, Z => snake_list(11));
  FE_OFC164_snake_list_7 : BUFFD5BWP7T port map(I => FE_OFN164_snake_list_7, Z => snake_list(7));
  FE_OFC163_snake_list_12 : BUFFD5BWP7T port map(I => FE_OFN163_snake_list_12, Z => snake_list(12));
  FE_OFC162_snake_list_9 : BUFFD5BWP7T port map(I => FE_OFN162_snake_list_9, Z => snake_list(9));
  FE_OFC161_snake_list_14 : BUFFD5BWP7T port map(I => FE_OFN161_snake_list_14, Z => snake_list(14));
  FE_OFC160_snake_list_6 : BUFFD5BWP7T port map(I => FE_OFN160_snake_list_6, Z => snake_list(6));
  FE_OFC159_snake_output24_5 : BUFFD5BWP7T port map(I => FE_OFN159_snake_output24_5, Z => snake_output24(5));
  FE_OFC158_snake_output24_1 : BUFFD5BWP7T port map(I => FE_OFN158_snake_output24_1, Z => snake_output24(1));
  FE_OFC157_snake_output24_2 : BUFFD5BWP7T port map(I => FE_OFN157_snake_output24_2, Z => snake_output24(2));
  FE_OFC156_snake_output24_4 : BUFFD5BWP7T port map(I => FE_OFN156_snake_output24_4, Z => snake_output24(4));
  FE_OFC155_snake_output24_0 : BUFFD5BWP7T port map(I => FE_OFN155_snake_output24_0, Z => snake_output24(0));
  FE_OFC154_snake_output24_3 : BUFFD5BWP7T port map(I => FE_OFN154_snake_output24_3, Z => snake_output24(3));
  FE_OFC153_snake_output3_5 : BUFFD5BWP7T port map(I => FE_OFN153_snake_output3_5, Z => snake_output3(5));
  FE_OFC152_snake_output6_5 : BUFFD5BWP7T port map(I => FE_OFN152_snake_output6_5, Z => snake_output6(5));
  FE_OFC151_snake_output22_5 : BUFFD5BWP7T port map(I => FE_OFN151_snake_output22_5, Z => snake_output22(5));
  FE_OFC150_snake_output7_5 : BUFFD5BWP7T port map(I => FE_OFN150_snake_output7_5, Z => snake_output7(5));
  FE_OFC149_snake_output5_5 : BUFFD5BWP7T port map(I => FE_OFN149_snake_output5_5, Z => snake_output5(5));
  FE_OFC148_snake_output2_5 : BUFFD5BWP7T port map(I => FE_OFN148_snake_output2_5, Z => snake_output2(5));
  FE_OFC147_snake_output21_5 : BUFFD5BWP7T port map(I => FE_OFN147_snake_output21_5, Z => snake_output21(5));
  FE_OFC146_snake_output20_5 : BUFFD5BWP7T port map(I => FE_OFN146_snake_output20_5, Z => snake_output20(5));
  FE_OFC145_snake_output15_5 : BUFFD5BWP7T port map(I => FE_OFN145_snake_output15_5, Z => snake_output15(5));
  FE_OFC144_snake_output9_5 : BUFFD5BWP7T port map(I => FE_OFN144_snake_output9_5, Z => snake_output9(5));
  FE_OFC143_snake_output10_5 : BUFFD5BWP7T port map(I => FE_OFN143_snake_output10_5, Z => snake_output10(5));
  FE_OFC142_snake_output14_5 : BUFFD6BWP7T port map(I => FE_OFN142_snake_output14_5, Z => snake_output14(5));
  FE_OFC141_snake_output18_5 : BUFFD5BWP7T port map(I => FE_OFN141_snake_output18_5, Z => snake_output18(5));
  FE_OFC140_snake_output12_5 : BUFFD5BWP7T port map(I => FE_OFN140_snake_output12_5, Z => snake_output12(5));
  FE_OFC139_snake_output13_5 : BUFFD6BWP7T port map(I => FE_OFN139_snake_output13_5, Z => snake_output13(5));
  FE_OFC138_snake_output19_5 : BUFFD6BWP7T port map(I => FE_OFN138_snake_output19_5, Z => snake_output19(5));
  FE_OFC137_snake_output16_5 : BUFFD6BWP7T port map(I => FE_OFN137_snake_output16_5, Z => snake_output16(5));
  FE_OFC136_snake_output17_5 : BUFFD6BWP7T port map(I => FE_OFN136_snake_output17_5, Z => snake_output17(5));
  FE_OFC135_snake_output11_5 : BUFFD6BWP7T port map(I => FE_OFN135_snake_output11_5, Z => snake_output11(5));
  FE_OFC134_snake_output8_5 : BUFFD6BWP7T port map(I => FE_OFN134_snake_output8_5, Z => snake_output8(5));
  FE_OFC133_snake_output23_0 : BUFFD5BWP7T port map(I => FE_OFN133_snake_output23_0, Z => snake_output23(0));
  FE_OFC132_snake_output23_3 : BUFFD5BWP7T port map(I => FE_OFN132_snake_output23_3, Z => snake_output23(3));
  FE_OFC131_snake_output23_1 : BUFFD5BWP7T port map(I => FE_OFN131_snake_output23_1, Z => snake_output23(1));
  FE_OFC130_snake_output23_4 : BUFFD5BWP7T port map(I => FE_OFN130_snake_output23_4, Z => snake_output23(4));
  FE_OFC129_snake_output21_3 : BUFFD5BWP7T port map(I => FE_OFN129_snake_output21_3, Z => snake_output21(3));
  FE_OFC128_snake_output23_2 : BUFFD5BWP7T port map(I => FE_OFN128_snake_output23_2, Z => snake_output23(2));
  FE_OFC127_snake_output20_3 : BUFFD5BWP7T port map(I => FE_OFN127_snake_output20_3, Z => snake_output20(3));
  FE_OFC126_snake_output20_1 : BUFFD5BWP7T port map(I => FE_OFN126_snake_output20_1, Z => snake_output20(1));
  FE_OFC125_snake_output22_1 : BUFFD5BWP7T port map(I => FE_OFN125_snake_output22_1, Z => snake_output22(1));
  FE_OFC124_snake_output20_0 : BUFFD5BWP7T port map(I => FE_OFN124_snake_output20_0, Z => snake_output20(0));
  FE_OFC123_snake_output19_1 : BUFFD5BWP7T port map(I => FE_OFN123_snake_output19_1, Z => snake_output19(1));
  FE_OFC122_snake_output22_3 : BUFFD5BWP7T port map(I => FE_OFN122_snake_output22_3, Z => snake_output22(3));
  FE_OFC121_snake_output21_4 : BUFFD5BWP7T port map(I => FE_OFN121_snake_output21_4, Z => snake_output21(4));
  FE_OFC120_snake_output21_1 : BUFFD5BWP7T port map(I => FE_OFN120_snake_output21_1, Z => snake_output21(1));
  FE_OFC119_snake_output20_4 : BUFFD5BWP7T port map(I => FE_OFN119_snake_output20_4, Z => snake_output20(4));
  FE_OFC118_snake_output22_0 : BUFFD5BWP7T port map(I => FE_OFN118_snake_output22_0, Z => snake_output22(0));
  FE_OFC117_snake_output22_4 : BUFFD5BWP7T port map(I => FE_OFN117_snake_output22_4, Z => snake_output22(4));
  FE_OFC116_snake_output18_1 : BUFFD5BWP7T port map(I => FE_OFN116_snake_output18_1, Z => snake_output18(1));
  FE_OFC115_snake_output18_4 : BUFFD5BWP7T port map(I => FE_OFN115_snake_output18_4, Z => snake_output18(4));
  FE_OFC114_snake_output1_2 : BUFFD5BWP7T port map(I => FE_OFN114_snake_output1_2, Z => snake_output1(2));
  FE_OFC113_snake_output1_3 : BUFFD5BWP7T port map(I => FE_OFN113_snake_output1_3, Z => snake_output1(3));
  FE_OFC112_snake_output19_3 : BUFFD5BWP7T port map(I => FE_OFN112_snake_output19_3, Z => snake_output19(3));
  FE_OFC111_snake_output19_4 : BUFFD5BWP7T port map(I => FE_OFN111_snake_output19_4, Z => snake_output19(4));
  FE_OFC110_snake_output20_2 : BUFFD5BWP7T port map(I => FE_OFN110_snake_output20_2, Z => snake_output20(2));
  FE_OFC109_snake_output2_2 : BUFFD5BWP7T port map(I => FE_OFN109_snake_output2_2, Z => snake_output2(2));
  FE_OFC108_snake_output17_4 : BUFFD5BWP7T port map(I => FE_OFN108_snake_output17_4, Z => snake_output17(4));
  FE_OFC107_snake_output17_3 : BUFFD5BWP7T port map(I => FE_OFN107_snake_output17_3, Z => snake_output17(3));
  FE_OFC106_snake_output16_1 : BUFFD5BWP7T port map(I => FE_OFN106_snake_output16_1, Z => snake_output16(1));
  FE_OFC105_snake_output5_4 : BUFFD5BWP7T port map(I => FE_OFN105_snake_output5_4, Z => snake_output5(4));
  FE_OFC104_snake_output5_3 : BUFFD5BWP7T port map(I => FE_OFN104_snake_output5_3, Z => snake_output5(3));
  FE_OFC103_snake_output18_3 : BUFFD5BWP7T port map(I => FE_OFN103_snake_output18_3, Z => snake_output18(3));
  FE_OFC102_snake_output1_1 : BUFFD5BWP7T port map(I => FE_OFN102_snake_output1_1, Z => snake_output1(1));
  FE_OFC101_snake_output2_3 : BUFFD5BWP7T port map(I => FE_OFN101_snake_output2_3, Z => snake_output2(3));
  FE_OFC100_snake_output21_2 : BUFFD5BWP7T port map(I => FE_OFN100_snake_output21_2, Z => snake_output21(2));
  FE_OFC99_snake_output1_0 : BUFFD5BWP7T port map(I => FE_OFN99_snake_output1_0, Z => snake_output1(0));
  FE_OFC98_snake_output17_1 : BUFFD5BWP7T port map(I => FE_OFN98_snake_output17_1, Z => snake_output17(1));
  FE_OFC97_snake_output1_4 : BUFFD5BWP7T port map(I => FE_OFN97_snake_output1_4, Z => snake_output1(4));
  FE_OFC96_snake_output22_2 : BUFFD5BWP7T port map(I => FE_OFN96_snake_output22_2, Z => snake_output22(2));
  FE_OFC95_snake_output7_3 : BUFFD5BWP7T port map(I => FE_OFN95_snake_output7_3, Z => snake_output7(3));
  FE_OFC94_snake_output21_0 : BUFFD5BWP7T port map(I => FE_OFN94_snake_output21_0, Z => snake_output21(0));
  FE_OFC93_snake_output7_2 : BUFFD5BWP7T port map(I => FE_OFN93_snake_output7_2, Z => snake_output7(2));
  FE_OFC92_snake_output3_2 : BUFFD5BWP7T port map(I => FE_OFN92_snake_output3_2, Z => snake_output3(2));
  FE_OFC91_snake_output16_3 : BUFFD5BWP7T port map(I => FE_OFN91_snake_output16_3, Z => snake_output16(3));
  FE_OFC90_snake_output19_2 : BUFFD5BWP7T port map(I => FE_OFN90_snake_output19_2, Z => snake_output19(2));
  FE_OFC89_snake_output6_0 : BUFFD5BWP7T port map(I => FE_OFN89_snake_output6_0, Z => snake_output6(0));
  FE_OFC88_snake_output4_3 : BUFFD5BWP7T port map(I => FE_OFN88_snake_output4_3, Z => snake_output4(3));
  FE_OFC87_snake_output5_2 : BUFFD5BWP7T port map(I => FE_OFN87_snake_output5_2, Z => snake_output5(2));
  FE_OFC86_snake_output5_1 : BUFFD5BWP7T port map(I => FE_OFN86_snake_output5_1, Z => snake_output5(1));
  FE_OFC85_snake_output2_1 : BUFFD5BWP7T port map(I => FE_OFN85_snake_output2_1, Z => snake_output2(1));
  FE_OFC84_snake_output17_0 : BUFFD5BWP7T port map(I => FE_OFN84_snake_output17_0, Z => snake_output17(0));
  FE_OFC83_snake_output6_4 : BUFFD5BWP7T port map(I => FE_OFN83_snake_output6_4, Z => snake_output6(4));
  FE_OFC82_snake_output5_0 : BUFFD5BWP7T port map(I => FE_OFN82_snake_output5_0, Z => snake_output5(0));
  FE_OFC81_snake_output16_4 : BUFFD5BWP7T port map(I => FE_OFN81_snake_output16_4, Z => snake_output16(4));
  FE_OFC80_snake_output3_1 : BUFFD5BWP7T port map(I => FE_OFN80_snake_output3_1, Z => snake_output3(1));
  FE_OFC79_snake_output6_3 : BUFFD5BWP7T port map(I => FE_OFN79_snake_output6_3, Z => snake_output6(3));
  FE_OFC78_snake_output3_3 : BUFFD5BWP7T port map(I => FE_OFN78_snake_output3_3, Z => snake_output3(3));
  FE_OFC77_snake_output4_2 : BUFFD5BWP7T port map(I => FE_OFN77_snake_output4_2, Z => snake_output4(2));
  FE_OFC76_snake_output3_4 : BUFFD5BWP7T port map(I => FE_OFN76_snake_output3_4, Z => snake_output3(4));
  FE_OFC75_snake_output4_0 : BUFFD5BWP7T port map(I => FE_OFN75_snake_output4_0, Z => snake_output4(0));
  FE_OFC74_snake_output7_0 : BUFFD5BWP7T port map(I => FE_OFN74_snake_output7_0, Z => snake_output7(0));
  FE_OFC73_snake_output16_0 : BUFFD5BWP7T port map(I => FE_OFN73_snake_output16_0, Z => snake_output16(0));
  FE_OFC72_snake_output2_0 : BUFFD5BWP7T port map(I => FE_OFN72_snake_output2_0, Z => snake_output2(0));
  FE_OFC71_snake_output2_4 : BUFFD5BWP7T port map(I => FE_OFN71_snake_output2_4, Z => snake_output2(4));
  FE_OFC70_snake_output7_4 : BUFFD5BWP7T port map(I => FE_OFN70_snake_output7_4, Z => snake_output7(4));
  FE_OFC69_snake_output4_4 : BUFFD5BWP7T port map(I => FE_OFN69_snake_output4_4, Z => snake_output4(4));
  FE_OFC68_snake_output6_2 : BUFFD5BWP7T port map(I => FE_OFN68_snake_output6_2, Z => snake_output6(2));
  FE_OFC67_snake_output3_0 : BUFFD5BWP7T port map(I => FE_OFN67_snake_output3_0, Z => snake_output3(0));
  FE_OFC66_snake_output4_1 : BUFFD5BWP7T port map(I => FE_OFN66_snake_output4_1, Z => snake_output4(1));
  FE_OFC65_snake_output12_1 : BUFFD5BWP7T port map(I => FE_OFN65_snake_output12_1, Z => snake_output12(1));
  FE_OFC64_snake_output6_1 : BUFFD5BWP7T port map(I => FE_OFN64_snake_output6_1, Z => snake_output6(1));
  FE_OFC63_snake_output11_2 : BUFFD5BWP7T port map(I => FE_OFN63_snake_output11_2, Z => snake_output11(2));
  FE_OFC62_snake_output19_0 : BUFFD5BWP7T port map(I => FE_OFN62_snake_output19_0, Z => snake_output19(0));
  FE_OFC61_snake_output18_0 : BUFFD5BWP7T port map(I => FE_OFN61_snake_output18_0, Z => snake_output18(0));
  FE_OFC60_snake_output12_3 : BUFFD5BWP7T port map(I => FE_OFN60_snake_output12_3, Z => snake_output12(3));
  FE_OFC59_snake_output12_2 : BUFFD5BWP7T port map(I => FE_OFN59_snake_output12_2, Z => snake_output12(2));
  FE_OFC58_snake_output11_3 : BUFFD5BWP7T port map(I => FE_OFN58_snake_output11_3, Z => snake_output11(3));
  FE_OFC57_snake_output13_2 : BUFFD5BWP7T port map(I => FE_OFN57_snake_output13_2, Z => snake_output13(2));
  FE_OFC56_snake_output10_2 : BUFFD5BWP7T port map(I => FE_OFN56_snake_output10_2, Z => snake_output10(2));
  FE_OFC55_snake_output11_1 : BUFFD5BWP7T port map(I => FE_OFN55_snake_output11_1, Z => snake_output11(1));
  FE_OFC54_snake_output13_3 : BUFFD5BWP7T port map(I => FE_OFN54_snake_output13_3, Z => snake_output13(3));
  FE_OFC53_snake_output11_4 : BUFFD5BWP7T port map(I => FE_OFN53_snake_output11_4, Z => snake_output11(4));
  FE_OFC52_snake_output11_0 : BUFFD5BWP7T port map(I => FE_OFN52_snake_output11_0, Z => snake_output11(0));
  FE_OFC51_snake_output18_2 : BUFFD5BWP7T port map(I => FE_OFN51_snake_output18_2, Z => snake_output18(2));
  FE_OFC50_snake_output15_1 : BUFFD5BWP7T port map(I => FE_OFN50_snake_output15_1, Z => snake_output15(1));
  FE_OFC49_snake_output15_2 : BUFFD5BWP7T port map(I => FE_OFN49_snake_output15_2, Z => snake_output15(2));
  FE_OFC48_snake_output10_4 : BUFFD5BWP7T port map(I => FE_OFN48_snake_output10_4, Z => snake_output10(4));
  FE_OFC47_snake_output13_1 : BUFFD5BWP7T port map(I => FE_OFN47_snake_output13_1, Z => snake_output13(1));
  FE_OFC46_snake_output17_2 : BUFFD5BWP7T port map(I => FE_OFN46_snake_output17_2, Z => snake_output17(2));
  FE_OFC45_snake_output9_3 : BUFFD5BWP7T port map(I => FE_OFN45_snake_output9_3, Z => snake_output9(3));
  FE_OFC44_snake_output7_1 : BUFFD5BWP7T port map(I => FE_OFN44_snake_output7_1, Z => snake_output7(1));
  FE_OFC43_snake_output9_4 : BUFFD5BWP7T port map(I => FE_OFN43_snake_output9_4, Z => snake_output9(4));
  FE_OFC42_snake_output10_0 : BUFFD5BWP7T port map(I => FE_OFN42_snake_output10_0, Z => snake_output10(0));
  FE_OFC41_snake_output16_2 : BUFFD5BWP7T port map(I => FE_OFN41_snake_output16_2, Z => snake_output16(2));
  FE_OFC40_snake_output12_4 : BUFFD5BWP7T port map(I => FE_OFN40_snake_output12_4, Z => snake_output12(4));
  FE_OFC39_snake_output15_3 : BUFFD5BWP7T port map(I => FE_OFN39_snake_output15_3, Z => snake_output15(3));
  FE_OFC38_snake_output13_4 : BUFFD5BWP7T port map(I => FE_OFN38_snake_output13_4, Z => snake_output13(4));
  FE_OFC37_snake_output13_0 : BUFFD5BWP7T port map(I => FE_OFN37_snake_output13_0, Z => snake_output13(0));
  FE_OFC36_snake_output9_1 : BUFFD5BWP7T port map(I => FE_OFN36_snake_output9_1, Z => snake_output9(1));
  FE_OFC35_snake_output9_2 : BUFFD5BWP7T port map(I => FE_OFN35_snake_output9_2, Z => snake_output9(2));
  FE_OFC34_snake_output14_1 : BUFFD5BWP7T port map(I => FE_OFN34_snake_output14_1, Z => snake_output14(1));
  FE_OFC33_snake_output1_5 : BUFFD5BWP7T port map(I => FE_OFN33_snake_output1_5, Z => snake_output1(5));
  FE_OFC32_snake_output14_2 : BUFFD5BWP7T port map(I => FE_OFN32_snake_output14_2, Z => snake_output14(2));
  FE_OFC31_snake_output12_0 : BUFFD5BWP7T port map(I => FE_OFN31_snake_output12_0, Z => snake_output12(0));
  FE_OFC30_snake_output10_3 : BUFFD6BWP7T port map(I => FE_OFN30_snake_output10_3, Z => snake_output10(3));
  FE_OFC29_snake_output10_1 : BUFFD6BWP7T port map(I => FE_OFN29_snake_output10_1, Z => snake_output10(1));
  FE_OFC28_snake_output14_4 : BUFFD5BWP7T port map(I => FE_OFN28_snake_output14_4, Z => snake_output14(4));
  FE_OFC27_snake_output14_0 : BUFFD5BWP7T port map(I => FE_OFN27_snake_output14_0, Z => snake_output14(0));
  FE_OFC26_snake_output9_0 : BUFFD5BWP7T port map(I => FE_OFN26_snake_output9_0, Z => snake_output9(0));
  FE_OFC25_snake_output8_3 : BUFFD5BWP7T port map(I => FE_OFN25_snake_output8_3, Z => snake_output8(3));
  FE_OFC24_snake_output15_4 : BUFFD5BWP7T port map(I => FE_OFN24_snake_output15_4, Z => snake_output15(4));
  FE_OFC23_snake_output14_3 : BUFFD5BWP7T port map(I => FE_OFN23_snake_output14_3, Z => snake_output14(3));
  FE_OFC22_snake_output15_0 : BUFFD5BWP7T port map(I => FE_OFN22_snake_output15_0, Z => snake_output15(0));
  FE_OFC21_snake_output8_4 : BUFFD5BWP7T port map(I => FE_OFN21_snake_output8_4, Z => snake_output8(4));
  FE_OFC20_snake_output8_0 : BUFFD5BWP7T port map(I => FE_OFN20_snake_output8_0, Z => snake_output8(0));
  FE_OFC19_snake_output8_1 : BUFFD5BWP7T port map(I => FE_OFN19_snake_output8_1, Z => snake_output8(1));
  FE_OFC18_snake_output8_2 : BUFFD5BWP7T port map(I => FE_OFN18_snake_output8_2, Z => snake_output8(2));
  FE_OFC17_audio_0 : BUFFD5BWP7T port map(I => audio(6), Z => audio(7));
  FE_OFC16_audio_0 : BUFFD5BWP7T port map(I => audio(5), Z => audio(6));
  FE_OFC15_audio_0 : BUFFD5BWP7T port map(I => audio(4), Z => audio(5));
  FE_OFC14_audio_0 : BUFFD5BWP7T port map(I => audio(3), Z => audio(4));
  FE_OFC13_audio_0 : BUFFD5BWP7T port map(I => item_send_flag, Z => send_new_corner_clear);
  FE_OFC12_audio_0 : BUFFD5BWP7T port map(I => audio(2), Z => audio(3));
  FE_OFC11_audio_0 : BUFFD5BWP7T port map(I => head_send_flag, Z => item_send_flag);
  FE_OFC10_audio_0 : BUFFD5BWP7T port map(I => audio(1), Z => audio(2));
  FE_OFC9_audio_0 : BUFFD5BWP7T port map(I => remove_item_clear, Z => head_send_flag);
  FE_OFC8_audio_0 : BUFFD5BWP7T port map(I => audio(0), Z => audio(1));
  FE_OFC7_audio_0 : INVD5BWP7T port map(I => FE_OFN6_audio_0, ZN => remove_item_clear);
  FE_OFC6_audio_0 : INVD5BWP7T port map(I => FE_OFN6_audio_0, ZN => FE_RN_11);
  FE_OFC5_audio_0 : INVD1BWP7T port map(I => FE_OFN5_audio_0, ZN => FE_OFN6_audio_0);
  FE_OFC4_n_1704 : BUFFD1P5BWP7T port map(I => FE_OFN3_n_1704, Z => FE_OFN4_n_1704);
  FE_OFC3_n_1704 : BUFFD1P5BWP7T port map(I => n_1704, Z => FE_OFN3_n_1704);
  FE_OFC2_n_1651 : BUFFD1P5BWP7T port map(I => n_1651, Z => FE_OFN2_n_1651);
  FE_OFC1_n_1657 : BUFFD2BWP7T port map(I => FE_OFN0_n_1657, Z => FE_OFN1_n_1657);
  FE_OFC0_n_1657 : BUFFD2BWP7T port map(I => n_1657, Z => FE_OFN0_n_1657);
  CTS_ccl_a_BUF_clk_G0_L1_1 : CKBD6BWP7T port map(I => clk, Z => CTS_6);
  g7522 : INVD5BWP7T port map(I => FE_OFN2_n_1651, ZN => snake_send_flag);
  H_S_reg_0_0 : LHD1BWP7T port map(D => n_1312, E => n_1353, Q => UNCONNECTED, QN => n_1350);
  H_S_reg_0_1 : LHD1BWP7T port map(D => n_1311, E => n_1353, Q => UNCONNECTED0, QN => n_1346);
  H_S_reg_0_2 : LHD1BWP7T port map(D => n_1310, E => n_1353, Q => UNCONNECTED1, QN => n_1347);
  H_S_reg_0_3 : LHD1BWP7T port map(D => n_1309, E => n_1353, Q => UNCONNECTED2, QN => n_1354);
  H_S_reg_0_4 : LHD1BWP7T port map(D => n_1313, E => n_1353, Q => UNCONNECTED3, QN => n_1351);
  H_S_reg_0_5 : LHD1BWP7T port map(D => n_1315, E => n_1353, Q => UNCONNECTED4, QN => n_1352);
  H_S_reg_0_6 : LHD1BWP7T port map(D => n_1314, E => n_1353, Q => UNCONNECTED5, QN => n_1337);
  H_S_reg_0_7 : LHD1BWP7T port map(D => n_1291, E => n_1353, Q => UNCONNECTED6, QN => n_1343);
  H_S_reg_0_8 : LHD1BWP7T port map(D => n_1292, E => n_1353, Q => UNCONNECTED7, QN => n_1348);
  H_S_reg_0_9 : LHD1BWP7T port map(D => n_1317, E => n_1353, Q => UNCONNECTED8, QN => n_1344);
  H_S_reg_0_10 : LHD1BWP7T port map(D => n_1300, E => n_1353, Q => UNCONNECTED9, QN => n_1345);
  H_S_reg_0_11 : LHD1BWP7T port map(D => n_1293, E => n_1353, Q => UNCONNECTED10, QN => n_1349);
  I_S_reg_0_0 : LHD1BWP7T port map(D => n_1301, E => n_1386, Q => UNCONNECTED11, QN => n_1366);
  I_S_reg_0_1 : LHD1BWP7T port map(D => n_1299, E => n_1386, Q => UNCONNECTED12, QN => n_1370);
  I_S_reg_0_2 : LHD1BWP7T port map(D => n_1319, E => n_1386, Q => UNCONNECTED13, QN => n_1374);
  I_S_reg_0_3 : LHD1BWP7T port map(D => n_1298, E => n_1386, Q => UNCONNECTED14, QN => n_1376);
  I_S_reg_0_4 : LHD1BWP7T port map(D => n_1297, E => n_1386, Q => UNCONNECTED15, QN => n_1380);
  I_S_reg_0_5 : LHD1BWP7T port map(D => n_1296, E => n_1386, Q => UNCONNECTED16, QN => n_1388);
  I_S_reg_0_6 : LHD1BWP7T port map(D => n_1316, E => n_1386, Q => UNCONNECTED17, QN => n_1365);
  I_S_reg_0_7 : LHD1BWP7T port map(D => n_1295, E => n_1386, Q => UNCONNECTED18, QN => n_1371);
  I_S_reg_0_8 : LHD1BWP7T port map(D => n_1294, E => n_1386, Q => UNCONNECTED19, QN => n_1377);
  I_S_reg_0_9 : LHD1BWP7T port map(D => n_1302, E => n_1386, Q => UNCONNECTED20, QN => n_1382);
  I_S_reg_0_10 : LHD1BWP7T port map(D => n_1327, E => n_1386, Q => UNCONNECTED21, QN => n_1368);
  I_S_reg_0_11 : LHD1BWP7T port map(D => n_1330, E => n_1386, Q => UNCONNECTED22, QN => n_1385);
  I_S_reg_1_0 : LND1BWP7T port map(D => n_1331, EN => n_1384, Q => UNCONNECTED23, QN => n_1367);
  I_S_reg_1_1 : LND1BWP7T port map(D => n_1329, EN => n_1384, Q => UNCONNECTED24, QN => n_1369);
  I_S_reg_1_2 : LND1BWP7T port map(D => n_1328, EN => n_1384, Q => UNCONNECTED25, QN => n_1372);
  I_S_reg_1_3 : LND1BWP7T port map(D => n_1318, EN => n_1384, Q => UNCONNECTED26, QN => n_1373);
  I_S_reg_1_4 : LND1BWP7T port map(D => n_1326, EN => n_1384, Q => UNCONNECTED27, QN => n_1375);
  I_S_reg_1_5 : LND1BWP7T port map(D => n_1325, EN => n_1384, Q => UNCONNECTED28, QN => n_1378);
  I_S_reg_1_6 : LND1BWP7T port map(D => n_1324, EN => n_1384, Q => UNCONNECTED29, QN => n_1379);
  I_S_reg_1_7 : LND1BWP7T port map(D => n_1332, EN => n_1384, Q => UNCONNECTED30, QN => n_1381);
  I_S_reg_1_8 : LND1BWP7T port map(D => n_1323, EN => n_1384, Q => UNCONNECTED31, QN => n_1383);
  I_S_reg_1_9 : LND1BWP7T port map(D => n_1322, EN => n_1384, Q => UNCONNECTED32, QN => n_1387);
  I_S_reg_1_10 : LND1BWP7T port map(D => n_1321, EN => n_1384, Q => UNCONNECTED33, QN => n_1363);
  I_S_reg_1_11 : LND1BWP7T port map(D => n_1320, EN => n_1384, Q => UNCONNECTED34, QN => n_1364);
  S_S_reg_0_0 : LND1BWP7T port map(D => n_1341, EN => n_1401, Q => UNCONNECTED35, QN => n_1400);
  S_S_reg_0_1 : LND1BWP7T port map(D => n_1360, EN => n_1401, Q => UNCONNECTED36, QN => n_1395);
  S_S_reg_0_2 : LND1BWP7T port map(D => n_1359, EN => n_1401, Q => UNCONNECTED37, QN => n_155);
  S_S_reg_0_3 : LND1BWP7T port map(D => n_1358, EN => n_1401, Q => UNCONNECTED38, QN => n_1402);
  S_S_reg_0_4 : LND1BWP7T port map(D => n_1357, EN => n_1401, Q => UNCONNECTED39, QN => n_1394);
  S_S_reg_0_5 : LND1BWP7T port map(D => n_1335, EN => n_1401, Q => UNCONNECTED40, QN => n_1399);
  new_N_reg_0 : LNQD1BWP7T port map(D => n_152, EN => FE_OFN2_n_1651, Q => new_N(0));
  new_corner_count_reg_0 : LHQD1BWP7T port map(D => n_146, E => FE_OFN0_n_1657, Q => new_corner_count(0));
  new_state_reg_2 : LHQD1BWP7T port map(D => n_1415, E => n_1649, Q => new_state(2));
  new_state_reg_3 : LHQD1BWP7T port map(D => n_1414, E => n_1649, Q => new_state(3));
  new_state_reg_4 : LHQD1BWP7T port map(D => n_1420, E => n_1649, Q => new_state(4));
  snake_list_reg_0 : LHD1BWP7T port map(D => n_1411, E => n_1652, Q => UNCONNECTED41, QN => n_1417);
  tail_reg : LHD1BWP7T port map(D => n_1404, E => FE_OFN2_n_1651, Q => UNCONNECTED42, QN => n_1407);
  g12536 : IND4D0BWP7T port map(A1 => n_1569, B1 => n_1279, B2 => n_1307, B3 => n_1426, ZN => n_1649);
  g12537 : NR4D0BWP7T port map(A1 => n_1425, A2 => n_1410, A3 => n_1579, A4 => n_1734, ZN => n_1426);
  g12538 : AO21D0BWP7T port map(A1 => n_1274, A2 => n_1209, B => n_1571, Z => n_1425);
  g12539 : AN2D1BWP7T port map(A1 => n_1650, A2 => n_1654, Z => n_1571);
  g12540 : IND4D0BWP7T port map(A1 => corner_count(8), B1 => n_1212, B2 => corner_count(0), B3 => n_1424, ZN => n_1650);
  g12541 : INR4D0BWP7T port map(A1 => n_1423, B1 => corner_count(9), B2 => corner_count(12), B3 => corner_count(10), ZN => n_1424);
  g12542 : INR4D0BWP7T port map(A1 => n_1422, B1 => corner_count(13), B2 => corner_count(16), B3 => corner_count(14), ZN => n_1423);
  g12543 : INR4D0BWP7T port map(A1 => n_1421, B1 => corner_count(17), B2 => corner_count(20), B3 => corner_count(18), ZN => n_1422);
  g12544 : INR4D0BWP7T port map(A1 => n_1419, B1 => corner_count(21), B2 => corner_count(5), B3 => corner_count(4), ZN => n_1421);
  g12545 : AN4D1BWP7T port map(A1 => n_1418, A2 => n_1277, A3 => n_1279, A4 => n_1203, Z => n_1420);
  g12546 : INR4D0BWP7T port map(A1 => n_1416, B1 => corner_count(6), B2 => corner_count(7), B3 => corner_count(3), ZN => n_1419);
  g12547 : NR4D0BWP7T port map(A1 => n_1749, A2 => n_1303, A3 => new_item_clear, A4 => clear_corner_flag, ZN => n_1418);
  g12549 : INVD5BWP7T port map(I => n_1417, ZN => snake_list(0));
  g12550 : INR4D0BWP7T port map(A1 => n_1408, B1 => corner_count(11), B2 => corner_count(19), B3 => corner_count(15), ZN => n_1416);
  g12551 : IND3D0BWP7T port map(A1 => n_1733, B1 => n_1409, B2 => n_1342, ZN => n_1415);
  g12552 : OR4D0BWP7T port map(A1 => n_1406, A2 => n_1734, A3 => n_1303, A4 => n_1568, Z => n_1414);
  g12553 : ND2D0BWP7T port map(A1 => n_1413, A2 => n_1279, ZN => n_1652);
  g12554 : NR2D0BWP7T port map(A1 => n_1410, A2 => n_1654, ZN => n_1413);
  g12556 : INR2D0BWP7T port map(A1 => tail, B1 => FE_OFN2_n_1651, ZN => n_1411);
  g12557 : AOI211D0BWP7T port map(A1 => n_1572, A2 => n_1747, B => n_1334, C => n_1403, ZN => n_1409);
  g12558 : IND4D0BWP7T port map(A1 => n_1572, B1 => n_1222, B2 => n_1276, B3 => n_1396, ZN => n_1410);
  g12559 : INR4D0BWP7T port map(A1 => n_1393, B1 => corner_count(22), B2 => corner_count(24), B3 => corner_count(23), ZN => n_1408);
  g12561 : INVD5BWP7T port map(I => n_1407, ZN => tail);
  g12562 : IND2D0BWP7T port map(A1 => n_1567, B1 => n_1392, ZN => n_1406);
  g12563 : OA221D0BWP7T port map(A1 => n_1283, A2 => n_1573, B1 => n_1397, B2 => FE_OFN2_n_1651, C => n_1336, Z => n_1405);
  g12564 : AN2D1BWP7T port map(A1 => n_1737, A2 => n_1397, Z => n_1566);
  g12565 : AN2D1BWP7T port map(A1 => n_1653, A2 => n_1397, Z => n_1567);
  g12566 : IAO21D0BWP7T port map(A1 => n_1569, A2 => n_1733, B => n_1397, ZN => n_1404);
  g12567 : OA21D0BWP7T port map(A1 => n_1737, A2 => n_1732, B => n_1397, Z => n_1403);
  g12569 : INVD5BWP7T port map(I => n_1402, ZN => snake_output0(3));
  g12571 : INVD5BWP7T port map(I => n_1400, ZN => snake_output0(0));
  g12573 : INVD5BWP7T port map(I => n_1399, ZN => snake_output0(5));
  g12575 : INVD5BWP7T port map(I => n_155, ZN => snake_output0(2));
  g12576 : NR4D0BWP7T port map(A1 => n_1391, A2 => n_1568, A3 => n_1303, A4 => n_1305, ZN => n_1396);
  g12578 : INVD5BWP7T port map(I => n_1395, ZN => snake_output0(1));
  g12580 : INVD5BWP7T port map(I => n_1394, ZN => snake_output0(4));
  g12581 : ND4D0BWP7T port map(A1 => n_1389, A2 => n_1390, A3 => n_1262, A4 => n_1215, ZN => n_1397);
  g12582 : NR4D0BWP7T port map(A1 => n_1361, A2 => corner_count(26), A3 => corner_count(25), A4 => corner_count(27), ZN => n_1393);
  g12583 : AOI32D0BWP7T port map(A1 => n_1572, A2 => n_1585, A3 => n_1273, B1 => n_1306, B2 => send_corner_flag, ZN => n_1392);
  g12584 : AOI211D0BWP7T port map(A1 => n_1362, A2 => n_1305, B => n_1278, C => n_1739, ZN => n_1401);
  g12585 : IIND4D0BWP7T port map(A1 => n_1663, A2 => new_item_clear, B1 => n_1287, B2 => n_1275, ZN => n_1391);
  g12586 : NR4D0BWP7T port map(A1 => n_1355, A2 => n_1284, A3 => n_1246, A4 => n_1244, ZN => n_1390);
  g12587 : NR4D0BWP7T port map(A1 => n_1338, A2 => n_1285, A3 => n_1289, A4 => n_1249, ZN => n_1389);
  g12589 : INVD5BWP7T port map(I => n_1388, ZN => item_out_food(5));
  g12591 : INVD5BWP7T port map(I => n_1387, ZN => item_out_power_up(9));
  g12593 : INVD5BWP7T port map(I => n_1385, ZN => item_out_food(11));
  g12595 : INVD5BWP7T port map(I => n_1383, ZN => item_out_power_up(8));
  g12597 : INVD5BWP7T port map(I => n_1382, ZN => item_out_food(9));
  g12599 : INVD5BWP7T port map(I => n_1381, ZN => item_out_power_up(7));
  g12601 : INVD5BWP7T port map(I => n_1380, ZN => item_out_food(4));
  g12603 : INVD5BWP7T port map(I => n_1379, ZN => item_out_power_up(6));
  g12605 : INVD5BWP7T port map(I => n_1378, ZN => item_out_power_up(5));
  g12607 : INVD5BWP7T port map(I => n_1377, ZN => item_out_food(8));
  g12609 : INVD5BWP7T port map(I => n_1376, ZN => item_out_food(3));
  g12611 : INVD5BWP7T port map(I => n_1375, ZN => item_out_power_up(4));
  g12613 : INVD5BWP7T port map(I => n_1374, ZN => item_out_food(2));
  g12615 : INVD5BWP7T port map(I => n_1373, ZN => item_out_power_up(3));
  g12617 : INVD5BWP7T port map(I => n_1372, ZN => item_out_power_up(2));
  g12619 : INVD5BWP7T port map(I => n_1371, ZN => item_out_food(7));
  g12621 : INVD5BWP7T port map(I => n_1370, ZN => item_out_food(1));
  g12623 : INVD5BWP7T port map(I => n_1369, ZN => item_out_power_up(1));
  g12625 : INVD5BWP7T port map(I => n_1368, ZN => item_out_food(10));
  g12627 : INVD5BWP7T port map(I => n_1367, ZN => item_out_power_up(0));
  g12629 : INVD5BWP7T port map(I => n_1366, ZN => item_out_food(0));
  g12631 : INVD5BWP7T port map(I => n_1365, ZN => item_out_food(6));
  g12633 : INVD5BWP7T port map(I => n_1364, ZN => item_out_power_up(11));
  g12635 : INVD5BWP7T port map(I => n_1363, ZN => item_out_power_up(10));
  g12636 : INR2D0BWP7T port map(A1 => n_1580, B1 => n_1339, ZN => n_1362);
  g12637 : IND2D0BWP7T port map(A1 => corner_count(28), B1 => n_1340, ZN => n_1361);
  g12638 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(1), B1 => n_1670, B2 => new_tail(1), C => n_1739, Z => n_1360);
  g12639 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(2), B1 => n_1670, B2 => new_tail(2), C => n_1739, Z => n_1359);
  g12640 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(3), B1 => n_1670, B2 => new_tail(3), C => n_1739, Z => n_1358);
  g12641 : AO221D0BWP7T port map(A1 => n_1278, A2 => new_corner(4), B1 => n_1670, B2 => new_tail(4), C => n_1739, Z => n_1357);
  g12643 : ND4D0BWP7T port map(A1 => n_1288, A2 => n_1290, A3 => n_1234, A4 => n_1233, ZN => n_1355);
  g12644 : IND3D0BWP7T port map(A1 => new_item_set, B1 => n_1211, B2 => n_1333, ZN => n_1585);
  g12647 : INVD5BWP7T port map(I => n_1354, ZN => head(3));
  g12649 : INVD5BWP7T port map(I => n_1352, ZN => head(5));
  g12651 : INVD5BWP7T port map(I => n_1351, ZN => head(4));
  g12653 : INVD5BWP7T port map(I => n_1350, ZN => head(0));
  g12655 : INVD5BWP7T port map(I => n_1349, ZN => head(11));
  g12657 : INVD5BWP7T port map(I => n_1348, ZN => head(8));
  g12660 : INVD5BWP7T port map(I => n_1347, ZN => head(2));
  g12662 : INVD5BWP7T port map(I => n_1346, ZN => head(1));
  g12664 : INVD5BWP7T port map(I => n_1345, ZN => head(10));
  g12666 : INVD5BWP7T port map(I => n_1344, ZN => head(9));
  g12668 : INVD5BWP7T port map(I => n_1343, ZN => head(7));
  g12669 : MOAI22D0BWP7T port map(A1 => n_1277, A2 => n_1209, B1 => n_1278, B2 => new_corner(0), ZN => n_1341);
  g12670 : ND2D5BWP7T port map(A1 => n_1304, A2 => n_1279, ZN => clear_tail_flag);
  g12671 : INR4D0BWP7T port map(A1 => n_1740, B1 => corner_count(29), B2 => corner_count(31), B3 => corner_count(30), ZN => n_1340);
  g12672 : OR4D0BWP7T port map(A1 => n_1581, A2 => n_1582, A3 => n_1583, A4 => n_1584, Z => n_1339);
  g12673 : ND4D0BWP7T port map(A1 => n_1286, A2 => n_1252, A3 => n_1240, A4 => n_1250, ZN => n_1338);
  g12675 : INVD5BWP7T port map(I => n_1337, ZN => head(6));
  g12676 : OAI21D0BWP7T port map(A1 => n_1280, A2 => n_1266, B => n_1225, ZN => n_1336);
  g12677 : AO22D0BWP7T port map(A1 => n_1278, A2 => new_corner(5), B1 => new_tail(5), B2 => n_1670, Z => n_1335);
  g12678 : NR2D0BWP7T port map(A1 => n_1307, A2 => send_corner_flag, ZN => n_1334);
  g12679 : AOI21D0BWP7T port map(A1 => n_1570, A2 => n_1217, B => n_1568, ZN => n_1342);
  g12680 : IND3D0BWP7T port map(A1 => n_1718, B1 => n_1276, B2 => n_1282, ZN => n_1386);
  g12681 : AOI211D1BWP7T port map(A1 => n_1264, A2 => n_1578, B => n_1705, C => n_1739, ZN => n_1384);
  g12683 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(7), Z => n_1332);
  g12684 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(0), Z => n_1331);
  g12685 : INR2D0BWP7T port map(A1 => new_item(11), B1 => n_1282, ZN => n_1330);
  g12686 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(1), Z => n_1329);
  g12687 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(2), Z => n_1328);
  g12688 : INR2D0BWP7T port map(A1 => new_item(10), B1 => n_1282, ZN => n_1327);
  g12689 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(4), Z => n_1326);
  g12690 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(5), Z => n_1325);
  g12691 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(6), Z => n_1324);
  g12692 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(8), Z => n_1323);
  g12693 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(9), Z => n_1322);
  g12694 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(10), Z => n_1321);
  g12695 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(11), Z => n_1320);
  g12696 : INR2D0BWP7T port map(A1 => new_item(2), B1 => n_1282, ZN => n_1319);
  g12698 : AN2D1BWP7T port map(A1 => n_1705, A2 => new_item(3), Z => n_1318);
  g12699 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(9), Z => n_1317);
  g12700 : INR2D0BWP7T port map(A1 => new_item(6), B1 => n_1282, ZN => n_1316);
  g12701 : IND2D0BWP7T port map(A1 => new_head(5), B1 => n_1731, ZN => n_1315);
  g12702 : INR2D0BWP7T port map(A1 => n_1736, B1 => n_1211, ZN => n_1564);
  g12703 : INR2D0BWP7T port map(A1 => n_1662, B1 => n_1211, ZN => n_1565);
  g12704 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(6), Z => n_1314);
  g12705 : IND2D0BWP7T port map(A1 => new_head(4), B1 => n_1731, ZN => n_1313);
  g12706 : IND2D0BWP7T port map(A1 => new_head(0), B1 => n_1731, ZN => n_1312);
  g12707 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(1), Z => n_1311);
  g12708 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(2), Z => n_1310);
  g12709 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(3), Z => n_1309);
  g12710 : AN2D1BWP7T port map(A1 => n_1273, A2 => new_item_set, Z => n_1574);
  g12711 : INR2D0BWP7T port map(A1 => n_1273, B1 => remove_item_set, ZN => n_1333);
  g12712 : CKND1BWP7T port map(I => n_1307, ZN => n_1306);
  g12713 : INVD1BWP7T port map(I => n_1305, ZN => n_1304);
  g12714 : INR2D0BWP7T port map(A1 => new_item(9), B1 => n_1282, ZN => n_1302);
  g12715 : INR2D0BWP7T port map(A1 => new_item(0), B1 => n_1282, ZN => n_1301);
  g12716 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(10), Z => n_1300);
  g12717 : INR2D0BWP7T port map(A1 => new_item(1), B1 => n_1282, ZN => n_1299);
  g12718 : INR2D0BWP7T port map(A1 => new_item(3), B1 => n_1282, ZN => n_1298);
  g12719 : INR2D0BWP7T port map(A1 => new_item(4), B1 => n_1282, ZN => n_1297);
  g12720 : INR2D0BWP7T port map(A1 => new_item(5), B1 => n_1282, ZN => n_1296);
  g12721 : INR2D0BWP7T port map(A1 => new_item(7), B1 => n_1282, ZN => n_1295);
  g12722 : INR2D0BWP7T port map(A1 => new_item(8), B1 => n_1282, ZN => n_1294);
  g12723 : IND2D0BWP7T port map(A1 => new_head(11), B1 => n_1731, ZN => n_1293);
  g12724 : IND2D0BWP7T port map(A1 => new_head(8), B1 => n_1731, ZN => n_1292);
  g12725 : AN2D1BWP7T port map(A1 => n_1731, A2 => new_head(7), Z => n_1291);
  g12726 : NR4D0BWP7T port map(A1 => n_1247, A2 => n_1248, A3 => n_1261, A4 => n_1251, ZN => n_1290);
  g12727 : ND4D0BWP7T port map(A1 => n_1231, A2 => n_1239, A3 => n_1258, A4 => n_1260, ZN => n_1289);
  g12728 : NR4D0BWP7T port map(A1 => n_1230, A2 => n_1232, A3 => n_1229, A4 => n_1257, ZN => n_1288);
  g12729 : OAI21D0BWP7T port map(A1 => n_1263, A2 => n_1264, B => n_1224, ZN => n_1287);
  g12730 : AOI211D0BWP7T port map(A1 => n_1207, A2 => N(4), B => n_1243, C => n_1259, ZN => n_1286);
  g12731 : ND4D0BWP7T port map(A1 => n_1235, A2 => n_1237, A3 => n_1242, A4 => n_1245, ZN => n_1285);
  g12732 : ND4D0BWP7T port map(A1 => n_1228, A2 => n_1241, A3 => n_1238, A4 => n_1236, ZN => n_1284);
  g12733 : AN4D1BWP7T port map(A1 => n_1255, A2 => n_1253, A3 => n_1254, A4 => n_1256, Z => n_1580);
  g12735 : OR2D0BWP7T port map(A1 => n_1732, A2 => n_1733, Z => n_1579);
  g12736 : ND2D0BWP7T port map(A1 => n_1280, A2 => n_1224, ZN => n_1307);
  g12737 : AOI21D0BWP7T port map(A1 => n_1267, A2 => n_1203, B => n_1216, ZN => n_1305);
  g12738 : OR2D0BWP7T port map(A1 => n_1704, A2 => n_1657, Z => n_1303);
  g12739 : OA21D0BWP7T port map(A1 => n_1263, A2 => n_1265, B => n_1225, Z => n_1569);
  g12740 : OR2D0BWP7T port map(A1 => n_1731, A2 => n_1278, Z => n_1568);
  g12741 : OAI221D0BWP7T port map(A1 => n_1227, A2 => n_1204, B1 => state(1), B2 => state(2), C => n_1224, ZN => n_1651);
  g12742 : ND2D0BWP7T port map(A1 => n_1281, A2 => n_1276, ZN => n_1353);
  g12743 : INVD1BWP7T port map(I => n_1283, ZN => n_1572);
  g12744 : INVD1BWP7T port map(I => n_1281, ZN => n_1731);
  g12745 : CKAN2D8BWP7T port map(A1 => n_1270, A2 => n_1578, Z => clear_head_flag);
  g12746 : AN2D1BWP7T port map(A1 => n_1265, A2 => n_1225, Z => n_1738);
  g12747 : INR2D0BWP7T port map(A1 => n_1264, B1 => n_1216, ZN => n_1663);
  g12748 : AN2D1BWP7T port map(A1 => n_1264, A2 => n_1224, Z => n_1653);
  g12749 : AN2D1BWP7T port map(A1 => n_1202, A2 => n_1273, Z => n_1575);
  g12750 : OR2D0BWP7T port map(A1 => n_1266, A2 => n_1264, Z => n_1570);
  g12751 : NR2XD1BWP7T port map(A1 => n_1203, A2 => n_1216, ZN => n_1703);
  g12752 : NR2D0BWP7T port map(A1 => n_1269, A2 => n_1226, ZN => n_1734);
  g12753 : AN2D1BWP7T port map(A1 => n_1266, A2 => n_1224, Z => n_1732);
  g12754 : INR2D0BWP7T port map(A1 => n_1266, B1 => n_1216, ZN => n_1654);
  g12756 : NR2D1P5BWP7T port map(A1 => n_1272, A2 => n_1216, ZN => n_1657);
  g12757 : AN2D1BWP7T port map(A1 => n_1264, A2 => n_1225, Z => n_1733);
  g12758 : ND2D0BWP7T port map(A1 => n_1265, A2 => n_1217, ZN => n_1283);
  g12759 : ND2D0BWP7T port map(A1 => n_1266, A2 => n_1578, ZN => n_1282);
  g12760 : ND2D0BWP7T port map(A1 => n_1263, A2 => n_1217, ZN => n_1281);
  g12761 : CKND1BWP7T port map(I => n_1670, ZN => n_1277);
  g12762 : INVD0BWP7T port map(I => n_1739, ZN => n_1276);
  g12763 : INR2D0BWP7T port map(A1 => n_1263, B1 => n_1226, ZN => n_1735);
  g12764 : OAI211D0BWP7T port map(A1 => state(3), A2 => n_1205, B => state(2), C => state(4), ZN => n_1275);
  g12765 : NR4D0BWP7T port map(A1 => new_tail(4), A2 => new_tail(3), A3 => new_tail(2), A4 => new_tail(1), ZN => n_1274);
  g12766 : NR2D0BWP7T port map(A1 => n_1267, A2 => n_1223, ZN => n_1662);
  g12767 : INR2D0BWP7T port map(A1 => n_1263, B1 => n_1222, ZN => n_1718);
  g12768 : ND2D0BWP7T port map(A1 => n_1267, A2 => n_1272, ZN => n_1280);
  g12769 : AN2D1BWP7T port map(A1 => n_1268, A2 => n_1578, Z => n_1704);
  g12770 : NR2D0BWP7T port map(A1 => n_1272, A2 => n_1223, ZN => n_1736);
  g12771 : OR4D0BWP7T port map(A1 => n_146, A2 => n_1701, A3 => n_1700, A4 => n_1699, Z => n_1581);
  g12772 : CKAN2D8BWP7T port map(A1 => n_1271, A2 => n_1578, Z => clear_corner_flag);
  g12773 : AN2D1BWP7T port map(A1 => n_1263, A2 => n_1224, Z => n_1737);
  g12774 : CKAN2D8BWP7T port map(A1 => n_1268, A2 => n_1224, Z => new_item_clear);
  g12775 : ND2D1BWP7T port map(A1 => n_1265, A2 => n_1224, ZN => n_1279);
  g12776 : INR2D0BWP7T port map(A1 => n_1265, B1 => n_1222, ZN => n_1278);
  g12777 : NR2XD0BWP7T port map(A1 => n_1267, A2 => n_1216, ZN => n_1670);
  g12778 : NR2D2P5BWP7T port map(A1 => n_1269, A2 => n_1216, ZN => n_1739);
  g12779 : NR2D1BWP7T port map(A1 => n_1267, A2 => n_1222, ZN => n_1705);
  g12780 : INVD0BWP7T port map(I => n_1271, ZN => n_1272);
  g12781 : INVD0BWP7T port map(I => n_1203, ZN => n_1270);
  g12782 : INVD1BWP7T port map(I => n_1269, ZN => n_1268);
  g12783 : MAOI22D0BWP7T port map(A1 => n_1214, A2 => N(5), B1 => n_1207, B2 => N(4), ZN => n_1262);
  g12784 : CKXOR2D0BWP7T port map(A1 => N(14), A2 => corner_count(14), Z => n_1261);
  g12785 : XNR2D1BWP7T port map(A1 => corner_count(8), A2 => N(8), ZN => n_1260);
  g12786 : CKXOR2D0BWP7T port map(A1 => N(29), A2 => corner_count(29), Z => n_1259);
  g12787 : XNR2D1BWP7T port map(A1 => corner_count(9), A2 => N(9), ZN => n_1258);
  g12788 : CKXOR2D0BWP7T port map(A1 => N(16), A2 => corner_count(16), Z => n_1257);
  g12789 : NR4D0BWP7T port map(A1 => n_1683, A2 => n_1684, A3 => n_1685, A4 => n_1686, ZN => n_1256);
  g12790 : NR4D0BWP7T port map(A1 => n_1671, A2 => n_1672, A3 => n_1673, A4 => n_1674, ZN => n_1255);
  g12791 : NR4D0BWP7T port map(A1 => n_1679, A2 => n_1680, A3 => n_1681, A4 => n_1682, ZN => n_1254);
  g12792 : NR4D0BWP7T port map(A1 => n_1675, A2 => n_1676, A3 => n_1677, A4 => n_1678, ZN => n_1253);
  g12793 : INR3D0BWP7T port map(A1 => remove_item_set, B1 => remove_item_type, B2 => new_item_set, ZN => n_1742);
  g12794 : AOI22D0BWP7T port map(A1 => corner_count(5), A2 => n_1208, B1 => n_1206, B2 => N(6), ZN => n_1252);
  g12795 : OR4D0BWP7T port map(A1 => n_1690, A2 => n_1689, A3 => n_1688, A4 => n_1687, Z => n_1584);
  g12796 : OR4D0BWP7T port map(A1 => n_1694, A2 => n_1693, A3 => n_1692, A4 => n_1691, Z => n_1583);
  g12797 : OR4D0BWP7T port map(A1 => n_1698, A2 => n_1697, A3 => n_1696, A4 => n_1695, Z => n_1582);
  g12799 : NR3D0BWP7T port map(A1 => new_head_flag, A2 => new_corner_flag, A3 => new_tail_flag, ZN => n_1273);
  g12800 : NR2XD0BWP7T port map(A1 => n_1221, A2 => n_1204, ZN => n_1271);
  g12802 : ND2D1BWP7T port map(A1 => n_1227, A2 => n_1204, ZN => n_1269);
  g12803 : ND2D1BWP7T port map(A1 => n_1218, A2 => state(2), ZN => n_1267);
  g12804 : INR2D0BWP7T port map(A1 => n_1227, B1 => n_1204, ZN => n_1266);
  g12805 : NR2XD0BWP7T port map(A1 => n_1219, A2 => state(2), ZN => n_1265);
  g12806 : NR2D0BWP7T port map(A1 => n_1221, A2 => state(2), ZN => n_1264);
  g12807 : NR2D0BWP7T port map(A1 => n_1220, A2 => state(2), ZN => n_1263);
  g12808 : CKXOR2D0BWP7T port map(A1 => N(12), A2 => corner_count(12), Z => n_1251);
  g12809 : XNR2D1BWP7T port map(A1 => corner_count(28), A2 => N(28), ZN => n_1250);
  g12810 : CKXOR2D0BWP7T port map(A1 => N(7), A2 => corner_count(7), Z => n_1249);
  g12811 : CKXOR2D0BWP7T port map(A1 => N(15), A2 => corner_count(15), Z => n_1248);
  g12812 : CKXOR2D0BWP7T port map(A1 => N(13), A2 => corner_count(13), Z => n_1247);
  g12813 : CKXOR2D0BWP7T port map(A1 => N(27), A2 => corner_count(27), Z => n_1246);
  g12814 : XNR2D1BWP7T port map(A1 => corner_count(3), A2 => N(3), ZN => n_1245);
  g12815 : CKXOR2D0BWP7T port map(A1 => N(25), A2 => corner_count(25), Z => n_1244);
  g12816 : CKXOR2D0BWP7T port map(A1 => N(31), A2 => corner_count(31), Z => n_1243);
  g12817 : XNR2D1BWP7T port map(A1 => corner_count(2), A2 => N(2), ZN => n_1242);
  g12818 : XNR2D1BWP7T port map(A1 => corner_count(21), A2 => N(21), ZN => n_1241);
  g12819 : XNR2D1BWP7T port map(A1 => corner_count(30), A2 => N(30), ZN => n_1240);
  g12820 : XNR2D1BWP7T port map(A1 => corner_count(10), A2 => N(10), ZN => n_1239);
  g12821 : XNR2D1BWP7T port map(A1 => corner_count(23), A2 => N(23), ZN => n_1238);
  g12822 : MAOI22D0BWP7T port map(A1 => n_1212, A2 => N(1), B1 => n_1212, B2 => N(1), ZN => n_1237);
  g12823 : XNR2D1BWP7T port map(A1 => corner_count(20), A2 => N(20), ZN => n_1236);
  g12824 : AOI22D0BWP7T port map(A1 => corner_count(0), A2 => n_152, B1 => n_146, B2 => N(0), ZN => n_1235);
  g12825 : XNR2D1BWP7T port map(A1 => corner_count(26), A2 => N(26), ZN => n_1234);
  g12826 : XNR2D1BWP7T port map(A1 => corner_count(24), A2 => N(24), ZN => n_1233);
  g12827 : CKXOR2D0BWP7T port map(A1 => N(19), A2 => corner_count(19), Z => n_1232);
  g12828 : XNR2D1BWP7T port map(A1 => corner_count(11), A2 => N(11), ZN => n_1231);
  g12829 : CKXOR2D0BWP7T port map(A1 => N(18), A2 => corner_count(18), Z => n_1230);
  g12830 : CKXOR2D0BWP7T port map(A1 => N(17), A2 => corner_count(17), Z => n_1229);
  g12831 : XNR2D1BWP7T port map(A1 => corner_count(22), A2 => N(22), ZN => n_1228);
  g12832 : MOAI22D0BWP7T port map(A1 => corner_count(1), A2 => corner_count(2), B1 => corner_count(1), B2 => corner_count(2), ZN => n_1740);
  g12833 : INVD0BWP7T port map(I => n_1226, ZN => n_1225);
  g12834 : INVD0BWP7T port map(I => n_1224, ZN => n_1223);
  g12835 : INVD0BWP7T port map(I => n_1578, ZN => n_1222);
  g12836 : NR2XD0BWP7T port map(A1 => state(0), A2 => state(1), ZN => n_1227);
  g12837 : ND2D0BWP7T port map(A1 => state(3), A2 => state(4), ZN => n_1226);
  g12838 : INR2XD0BWP7T port map(A1 => state(4), B1 => state(3), ZN => n_1224);
  g12839 : INR2XD0BWP7T port map(A1 => state(3), B1 => state(4), ZN => n_1578);
  g12841 : INVD0BWP7T port map(I => n_1218, ZN => n_1219);
  g12842 : INVD1BWP7T port map(I => n_1217, ZN => n_1216);
  g12843 : IND2D0BWP7T port map(A1 => N(6), B1 => corner_count(6), ZN => n_1215);
  g12844 : ND2D1BWP7T port map(A1 => state(1), A2 => state(0), ZN => n_1221);
  g12845 : ND2D1BWP7T port map(A1 => n_1205, A2 => state(1), ZN => n_1220);
  g12846 : NR2XD0BWP7T port map(A1 => n_1205, A2 => state(1), ZN => n_1218);
  g12847 : NR2XD0BWP7T port map(A1 => state(4), A2 => state(3), ZN => n_1217);
  g12848 : CKND1BWP7T port map(I => corner_count(5), ZN => n_1214);
  g12850 : INVD0BWP7T port map(I => corner_count(1), ZN => n_1212);
  g12853 : INVD1BWP7T port map(I => send_corner_flag, ZN => n_1211);
  g12854 : INVD0BWP7T port map(I => new_head_flag, ZN => n_1210);
  g12855 : CKND1BWP7T port map(I => new_tail(0), ZN => n_1209);
  g12856 : CKND1BWP7T port map(I => N(5), ZN => n_1208);
  g12857 : CKND1BWP7T port map(I => corner_count(4), ZN => n_1207);
  g12858 : CKND1BWP7T port map(I => corner_count(6), ZN => n_1206);
  g2 : INR3D0BWP7T port map(A1 => n_1333, B1 => new_item_set, B2 => n_1211, ZN => n_1573);
  g12861 : IND2D1BWP7T port map(A1 => n_1220, B1 => state(2), ZN => n_1203);
  g12862 : INR3D0BWP7T port map(A1 => new_item_set, B1 => new_item(0), B2 => new_item(1), ZN => n_1202);
  N_reg_0 : LNQD1BWP7T port map(D => n_190, EN => FE_OFN176_n_483, Q => N(0));
  N_reg_1 : LNQD1BWP7T port map(D => n_162, EN => FE_OFN176_n_483, Q => N(1));
  N_reg_2 : LNQD1BWP7T port map(D => n_163, EN => FE_OFN176_n_483, Q => N(2));
  N_reg_3 : LNQD1BWP7T port map(D => n_191, EN => FE_OFN176_n_483, Q => N(3));
  N_reg_4 : LNQD1BWP7T port map(D => n_165, EN => FE_OFN176_n_483, Q => N(4));
  N_reg_5 : LNQD1BWP7T port map(D => n_169, EN => FE_OFN176_n_483, Q => N(5));
  N_reg_6 : LNQD1BWP7T port map(D => n_170, EN => FE_OFN176_n_483, Q => N(6));
  N_reg_7 : LNQD1BWP7T port map(D => n_173, EN => FE_OFN176_n_483, Q => N(7));
  N_reg_8 : LNQD1BWP7T port map(D => n_160, EN => FE_OFN176_n_483, Q => N(8));
  N_reg_9 : LNQD1BWP7T port map(D => n_159, EN => FE_OFN176_n_483, Q => N(9));
  N_reg_10 : LNQD1BWP7T port map(D => n_174, EN => FE_OFN176_n_483, Q => N(10));
  N_reg_11 : LNQD1BWP7T port map(D => n_167, EN => FE_OFN176_n_483, Q => N(11));
  N_reg_12 : LNQD1BWP7T port map(D => n_172, EN => FE_OFN176_n_483, Q => N(12));
  N_reg_13 : LNQD1BWP7T port map(D => n_178, EN => FE_OFN176_n_483, Q => N(13));
  N_reg_14 : LNQD1BWP7T port map(D => n_175, EN => FE_OFN176_n_483, Q => N(14));
  N_reg_15 : LNQD1BWP7T port map(D => n_177, EN => FE_OFN176_n_483, Q => N(15));
  N_reg_16 : LNQD1BWP7T port map(D => n_180, EN => FE_OFN176_n_483, Q => N(16));
  N_reg_17 : LNQD1BWP7T port map(D => n_166, EN => FE_OFN176_n_483, Q => N(17));
  N_reg_18 : LNQD1BWP7T port map(D => n_176, EN => FE_OFN176_n_483, Q => N(18));
  N_reg_19 : LNQD1BWP7T port map(D => n_179, EN => FE_OFN176_n_483, Q => N(19));
  N_reg_20 : LNQD1BWP7T port map(D => n_181, EN => FE_OFN176_n_483, Q => N(20));
  N_reg_21 : LNQD1BWP7T port map(D => n_171, EN => FE_OFN176_n_483, Q => N(21));
  N_reg_22 : LNQD1BWP7T port map(D => n_161, EN => FE_OFN176_n_483, Q => N(22));
  N_reg_23 : LNQD1BWP7T port map(D => n_158, EN => FE_OFN176_n_483, Q => N(23));
  N_reg_24 : LNQD1BWP7T port map(D => n_183, EN => FE_OFN176_n_483, Q => N(24));
  N_reg_25 : LNQD1BWP7T port map(D => n_168, EN => FE_OFN176_n_483, Q => N(25));
  N_reg_26 : LNQD1BWP7T port map(D => n_184, EN => FE_OFN176_n_483, Q => N(26));
  N_reg_27 : LNQD1BWP7T port map(D => n_185, EN => FE_OFN176_n_483, Q => N(27));
  N_reg_28 : LNQD1BWP7T port map(D => n_186, EN => FE_OFN176_n_483, Q => N(28));
  N_reg_29 : LNQD1BWP7T port map(D => n_182, EN => FE_OFN176_n_483, Q => N(29));
  N_reg_30 : LNQD1BWP7T port map(D => n_188, EN => FE_OFN176_n_483, Q => N(30));
  N_reg_31 : LNQD1BWP7T port map(D => n_189, EN => FE_OFN176_n_483, Q => N(31));
  S_S_reg_1_0 : LHQD1BWP7T port map(D => n_279, E => FE_OFN177_n_674, Q => FE_OFN99_snake_output1_0);
  S_S_reg_1_1 : LHQD1BWP7T port map(D => n_393, E => FE_OFN177_n_674, Q => FE_OFN102_snake_output1_1);
  S_S_reg_1_2 : LHQD1BWP7T port map(D => n_388, E => FE_OFN177_n_674, Q => FE_OFN114_snake_output1_2);
  S_S_reg_1_3 : LHQD1BWP7T port map(D => n_386, E => FE_OFN177_n_674, Q => FE_OFN113_snake_output1_3);
  S_S_reg_1_4 : LHQD1BWP7T port map(D => n_381, E => FE_OFN177_n_674, Q => FE_OFN97_snake_output1_4);
  S_S_reg_1_5 : LHQD1BWP7T port map(D => n_374, E => FE_OFN177_n_674, Q => FE_OFN33_snake_output1_5);
  S_S_reg_2_0 : LHQD1BWP7T port map(D => n_376, E => n_764, Q => FE_OFN72_snake_output2_0);
  S_S_reg_2_1 : LHQD1BWP7T port map(D => n_348, E => n_764, Q => FE_OFN85_snake_output2_1);
  S_S_reg_2_2 : LHQD1BWP7T port map(D => n_370, E => n_764, Q => FE_OFN109_snake_output2_2);
  S_S_reg_2_3 : LHQD1BWP7T port map(D => n_367, E => n_764, Q => FE_OFN101_snake_output2_3);
  S_S_reg_2_4 : LHQD1BWP7T port map(D => n_363, E => n_764, Q => FE_OFN71_snake_output2_4);
  S_S_reg_2_5 : LHQD1BWP7T port map(D => n_410, E => n_764, Q => FE_OFN148_snake_output2_5);
  S_S_reg_3_0 : LHQD1BWP7T port map(D => n_396, E => n_766, Q => FE_OFN67_snake_output3_0);
  S_S_reg_3_1 : LHQD1BWP7T port map(D => n_353, E => n_766, Q => FE_OFN80_snake_output3_1);
  S_S_reg_3_2 : LHQD1BWP7T port map(D => n_355, E => n_766, Q => FE_OFN92_snake_output3_2);
  S_S_reg_3_3 : LHQD1BWP7T port map(D => n_294, E => n_766, Q => FE_OFN78_snake_output3_3);
  S_S_reg_3_4 : LHQD1BWP7T port map(D => n_352, E => n_766, Q => FE_OFN76_snake_output3_4);
  S_S_reg_3_5 : LHQD1BWP7T port map(D => n_350, E => n_766, Q => FE_OFN153_snake_output3_5);
  S_S_reg_4_0 : LNQD1BWP7T port map(D => n_349, EN => n_598, Q => FE_OFN75_snake_output4_0);
  S_S_reg_4_1 : LNQD1BWP7T port map(D => n_298, EN => n_598, Q => FE_OFN66_snake_output4_1);
  S_S_reg_4_2 : LNQD1BWP7T port map(D => n_345, EN => n_598, Q => FE_OFN77_snake_output4_2);
  S_S_reg_4_3 : LNQD1BWP7T port map(D => n_344, EN => n_598, Q => FE_OFN88_snake_output4_3);
  S_S_reg_4_4 : LNQD1BWP7T port map(D => n_343, EN => n_598, Q => FE_OFN69_snake_output4_4);
  S_S_reg_4_5 : LNQD1BWP7T port map(D => n_356, EN => n_598, Q => n_1167);
  S_S_reg_5_0 : LNQD1BWP7T port map(D => n_394, EN => n_673, Q => FE_OFN82_snake_output5_0);
  S_S_reg_5_1 : LNQD1BWP7T port map(D => n_401, EN => n_673, Q => FE_OFN86_snake_output5_1);
  S_S_reg_5_2 : LNQD1BWP7T port map(D => n_398, EN => n_673, Q => FE_OFN87_snake_output5_2);
  S_S_reg_5_3 : LNQD1BWP7T port map(D => n_335, EN => n_673, Q => FE_OFN104_snake_output5_3);
  S_S_reg_5_4 : LNQD1BWP7T port map(D => n_395, EN => n_673, Q => FE_OFN105_snake_output5_4);
  S_S_reg_5_5 : LNQD1BWP7T port map(D => n_375, EN => n_673, Q => FE_OFN149_snake_output5_5);
  S_S_reg_6_0 : LHQD1BWP7T port map(D => n_321, E => n_765, Q => FE_OFN89_snake_output6_0);
  S_S_reg_6_1 : LHQD1BWP7T port map(D => n_284, E => n_765, Q => FE_OFN64_snake_output6_1);
  S_S_reg_6_2 : LHQD1BWP7T port map(D => n_286, E => n_765, Q => FE_OFN68_snake_output6_2);
  S_S_reg_6_3 : LHQD1BWP7T port map(D => n_413, E => n_765, Q => FE_OFN79_snake_output6_3);
  S_S_reg_6_4 : LHQD1BWP7T port map(D => n_354, E => n_765, Q => FE_OFN83_snake_output6_4);
  S_S_reg_6_5 : LHQD1BWP7T port map(D => n_288, E => n_765, Q => FE_OFN152_snake_output6_5);
  S_S_reg_7_0 : LHQD1BWP7T port map(D => n_406, E => n_763, Q => FE_OFN74_snake_output7_0);
  S_S_reg_7_1 : LHQD1BWP7T port map(D => n_399, E => n_763, Q => FE_OFN44_snake_output7_1);
  S_S_reg_7_2 : LHQD1BWP7T port map(D => n_402, E => n_763, Q => FE_OFN93_snake_output7_2);
  S_S_reg_7_3 : LHQD1BWP7T port map(D => n_403, E => n_763, Q => FE_OFN95_snake_output7_3);
  S_S_reg_7_4 : LHQD1BWP7T port map(D => n_404, E => n_763, Q => FE_OFN70_snake_output7_4);
  S_S_reg_7_5 : LHQD1BWP7T port map(D => n_308, E => n_763, Q => FE_OFN150_snake_output7_5);
  S_S_reg_8_0 : LNQD1BWP7T port map(D => n_342, EN => n_762, Q => FE_OFN20_snake_output8_0);
  S_S_reg_8_1 : LNQD1BWP7T port map(D => n_405, EN => n_762, Q => FE_OFN19_snake_output8_1);
  S_S_reg_8_2 : LNQD1BWP7T port map(D => n_319, EN => n_762, Q => FE_OFN18_snake_output8_2);
  S_S_reg_8_3 : LNQD1BWP7T port map(D => n_408, EN => n_762, Q => FE_OFN25_snake_output8_3);
  S_S_reg_8_4 : LNQD1BWP7T port map(D => n_409, EN => n_762, Q => FE_OFN21_snake_output8_4);
  S_S_reg_8_5 : LNQD1BWP7T port map(D => n_411, EN => n_762, Q => FE_OFN134_snake_output8_5);
  S_S_reg_9_0 : LNQD1BWP7T port map(D => n_397, EN => n_761, Q => FE_OFN26_snake_output9_0);
  S_S_reg_9_1 : LNQD1BWP7T port map(D => n_412, EN => n_761, Q => FE_OFN36_snake_output9_1);
  S_S_reg_9_2 : LNQD1BWP7T port map(D => n_400, EN => n_761, Q => FE_OFN35_snake_output9_2);
  S_S_reg_9_3 : LNQD1BWP7T port map(D => n_414, EN => n_761, Q => FE_OFN45_snake_output9_3);
  S_S_reg_9_4 : LNQD1BWP7T port map(D => n_360, EN => n_761, Q => FE_OFN43_snake_output9_4);
  S_S_reg_9_5 : LNQD1BWP7T port map(D => n_415, EN => n_761, Q => FE_OFN144_snake_output9_5);
  S_S_reg_10_0 : LNQD1BWP7T port map(D => n_328, EN => n_760, Q => FE_OFN42_snake_output10_0);
  S_S_reg_10_1 : LNQD1BWP7T port map(D => n_416, EN => n_760, Q => FE_OFN29_snake_output10_1);
  S_S_reg_10_2 : LNQD1BWP7T port map(D => n_340, EN => n_760, Q => FE_OFN56_snake_output10_2);
  S_S_reg_10_3 : LNQD1BWP7T port map(D => n_339, EN => n_760, Q => FE_OFN30_snake_output10_3);
  S_S_reg_10_4 : LNQD1BWP7T port map(D => n_338, EN => n_760, Q => FE_OFN48_snake_output10_4);
  S_S_reg_10_5 : LNQD1BWP7T port map(D => n_337, EN => n_760, Q => FE_OFN143_snake_output10_5);
  S_S_reg_11_0 : LNQD1BWP7T port map(D => n_336, EN => n_759, Q => FE_OFN52_snake_output11_0);
  S_S_reg_11_1 : LNQD1BWP7T port map(D => n_334, EN => n_759, Q => FE_OFN55_snake_output11_1);
  S_S_reg_11_2 : LNQD1BWP7T port map(D => n_333, EN => n_759, Q => FE_OFN63_snake_output11_2);
  S_S_reg_11_3 : LNQD1BWP7T port map(D => n_332, EN => n_759, Q => FE_OFN58_snake_output11_3);
  S_S_reg_11_4 : LNQD1BWP7T port map(D => n_331, EN => n_759, Q => FE_OFN53_snake_output11_4);
  S_S_reg_11_5 : LNQD1BWP7T port map(D => n_330, EN => n_759, Q => FE_OFN135_snake_output11_5);
  S_S_reg_12_0 : LNQD1BWP7T port map(D => n_329, EN => n_758, Q => FE_OFN31_snake_output12_0);
  S_S_reg_12_1 : LNQD1BWP7T port map(D => n_327, EN => n_758, Q => FE_OFN65_snake_output12_1);
  S_S_reg_12_2 : LNQD1BWP7T port map(D => n_326, EN => n_758, Q => FE_OFN59_snake_output12_2);
  S_S_reg_12_3 : LNQD1BWP7T port map(D => n_325, EN => n_758, Q => FE_OFN60_snake_output12_3);
  S_S_reg_12_4 : LNQD1BWP7T port map(D => n_324, EN => n_758, Q => FE_OFN40_snake_output12_4);
  S_S_reg_12_5 : LNQD1BWP7T port map(D => n_323, EN => n_758, Q => FE_OFN140_snake_output12_5);
  S_S_reg_13_0 : LNQD1BWP7T port map(D => n_322, EN => n_757, Q => FE_OFN37_snake_output13_0);
  S_S_reg_13_1 : LNQD1BWP7T port map(D => n_320, EN => n_757, Q => FE_OFN47_snake_output13_1);
  S_S_reg_13_2 : LNQD1BWP7T port map(D => n_318, EN => n_757, Q => FE_OFN57_snake_output13_2);
  S_S_reg_13_3 : LNQD1BWP7T port map(D => n_317, EN => n_757, Q => FE_OFN54_snake_output13_3);
  S_S_reg_13_4 : LNQD1BWP7T port map(D => n_316, EN => n_757, Q => FE_OFN38_snake_output13_4);
  S_S_reg_13_5 : LNQD1BWP7T port map(D => n_315, EN => n_757, Q => FE_OFN139_snake_output13_5);
  S_S_reg_14_0 : LHQD1BWP7T port map(D => n_314, E => n_756, Q => FE_OFN27_snake_output14_0);
  S_S_reg_14_1 : LHQD1BWP7T port map(D => n_313, E => n_756, Q => FE_OFN34_snake_output14_1);
  S_S_reg_14_2 : LHQD1BWP7T port map(D => n_312, E => n_756, Q => FE_OFN32_snake_output14_2);
  S_S_reg_14_3 : LHQD1BWP7T port map(D => n_311, E => n_756, Q => FE_OFN23_snake_output14_3);
  S_S_reg_14_4 : LHQD1BWP7T port map(D => n_310, E => n_756, Q => FE_OFN28_snake_output14_4);
  S_S_reg_14_5 : LHQD1BWP7T port map(D => n_309, E => n_756, Q => FE_OFN142_snake_output14_5);
  S_S_reg_15_0 : LHQD1BWP7T port map(D => n_307, E => n_702, Q => FE_OFN22_snake_output15_0);
  S_S_reg_15_1 : LHQD1BWP7T port map(D => n_306, E => n_702, Q => FE_OFN50_snake_output15_1);
  S_S_reg_15_2 : LHQD1BWP7T port map(D => n_305, E => n_702, Q => FE_OFN49_snake_output15_2);
  S_S_reg_15_3 : LHQD1BWP7T port map(D => n_304, E => n_702, Q => FE_OFN39_snake_output15_3);
  S_S_reg_15_4 : LHQD1BWP7T port map(D => n_303, E => n_702, Q => FE_OFN24_snake_output15_4);
  S_S_reg_15_5 : LHQD1BWP7T port map(D => n_302, E => n_702, Q => FE_OFN145_snake_output15_5);
  S_S_reg_16_0 : LHQD1BWP7T port map(D => n_301, E => n_812, Q => FE_OFN73_snake_output16_0);
  S_S_reg_16_1 : LHQD1BWP7T port map(D => n_300, E => n_812, Q => FE_OFN106_snake_output16_1);
  S_S_reg_16_2 : LHQD1BWP7T port map(D => n_299, E => n_812, Q => FE_OFN41_snake_output16_2);
  S_S_reg_16_3 : LHQD1BWP7T port map(D => n_297, E => n_812, Q => FE_OFN91_snake_output16_3);
  S_S_reg_16_4 : LHQD1BWP7T port map(D => n_296, E => n_812, Q => FE_OFN81_snake_output16_4);
  S_S_reg_16_5 : LHQD1BWP7T port map(D => n_295, E => n_812, Q => FE_OFN137_snake_output16_5);
  S_S_reg_17_0 : LHQD1BWP7T port map(D => n_407, E => n_859, Q => FE_OFN84_snake_output17_0);
  S_S_reg_17_1 : LHQD1BWP7T port map(D => n_293, E => n_859, Q => FE_OFN98_snake_output17_1);
  S_S_reg_17_2 : LHQD1BWP7T port map(D => n_292, E => n_859, Q => FE_OFN46_snake_output17_2);
  S_S_reg_17_3 : LHQD1BWP7T port map(D => n_291, E => n_859, Q => FE_OFN107_snake_output17_3);
  S_S_reg_17_4 : LHQD1BWP7T port map(D => n_290, E => n_859, Q => FE_OFN108_snake_output17_4);
  S_S_reg_17_5 : LHQD1BWP7T port map(D => n_289, E => n_859, Q => FE_OFN136_snake_output17_5);
  S_S_reg_18_0 : LNQD1BWP7T port map(D => n_287, EN => n_887, Q => FE_OFN61_snake_output18_0);
  S_S_reg_18_1 : LNQD1BWP7T port map(D => n_285, EN => n_887, Q => FE_OFN116_snake_output18_1);
  S_S_reg_18_2 : LNQD1BWP7T port map(D => n_283, EN => n_887, Q => FE_OFN51_snake_output18_2);
  S_S_reg_18_3 : LNQD1BWP7T port map(D => n_282, EN => n_887, Q => FE_OFN103_snake_output18_3);
  S_S_reg_18_4 : LNQD1BWP7T port map(D => n_281, EN => n_887, Q => FE_OFN115_snake_output18_4);
  S_S_reg_18_5 : LNQD1BWP7T port map(D => n_280, EN => n_887, Q => FE_OFN141_snake_output18_5);
  S_S_reg_19_0 : LNQD1BWP7T port map(D => n_278, EN => n_886, Q => FE_OFN62_snake_output19_0);
  S_S_reg_19_1 : LNQD1BWP7T port map(D => n_277, EN => n_886, Q => FE_OFN123_snake_output19_1);
  S_S_reg_19_2 : LNQD1BWP7T port map(D => n_276, EN => n_886, Q => FE_OFN90_snake_output19_2);
  S_S_reg_19_3 : LNQD1BWP7T port map(D => n_275, EN => n_886, Q => FE_OFN112_snake_output19_3);
  S_S_reg_19_4 : LNQD1BWP7T port map(D => n_274, EN => n_886, Q => FE_OFN111_snake_output19_4);
  S_S_reg_19_5 : LNQD1BWP7T port map(D => n_273, EN => n_886, Q => FE_OFN138_snake_output19_5);
  S_S_reg_20_0 : LHQD1BWP7T port map(D => n_392, E => n_811, Q => FE_OFN124_snake_output20_0);
  S_S_reg_20_1 : LHQD1BWP7T port map(D => n_391, E => n_811, Q => FE_OFN126_snake_output20_1);
  S_S_reg_20_2 : LHQD1BWP7T port map(D => n_390, E => n_811, Q => FE_OFN110_snake_output20_2);
  S_S_reg_20_3 : LHQD1BWP7T port map(D => n_389, E => n_811, Q => FE_OFN127_snake_output20_3);
  S_S_reg_20_4 : LHQD1BWP7T port map(D => n_387, E => n_811, Q => FE_OFN119_snake_output20_4);
  S_S_reg_20_5 : LHQD1BWP7T port map(D => n_385, E => n_811, Q => FE_OFN146_snake_output20_5);
  S_S_reg_21_0 : LNQD1BWP7T port map(D => n_384, EN => n_860, Q => FE_OFN94_snake_output21_0);
  S_S_reg_21_1 : LNQD1BWP7T port map(D => n_383, EN => n_860, Q => FE_OFN120_snake_output21_1);
  S_S_reg_21_2 : LNQD1BWP7T port map(D => n_382, EN => n_860, Q => FE_OFN100_snake_output21_2);
  S_S_reg_21_3 : LNQD1BWP7T port map(D => n_380, EN => n_860, Q => FE_OFN129_snake_output21_3);
  S_S_reg_21_4 : LNQD1BWP7T port map(D => n_379, EN => n_860, Q => FE_OFN121_snake_output21_4);
  S_S_reg_21_5 : LNQD1BWP7T port map(D => n_378, EN => n_860, Q => FE_OFN147_snake_output21_5);
  S_S_reg_22_0 : LHQD1BWP7T port map(D => n_377, E => n_889, Q => FE_OFN118_snake_output22_0);
  S_S_reg_22_1 : LHQD1BWP7T port map(D => n_373, E => n_889, Q => FE_OFN125_snake_output22_1);
  S_S_reg_22_2 : LHQD1BWP7T port map(D => n_372, E => n_889, Q => FE_OFN96_snake_output22_2);
  S_S_reg_22_3 : LHQD1BWP7T port map(D => n_371, E => n_889, Q => FE_OFN122_snake_output22_3);
  S_S_reg_22_4 : LHQD1BWP7T port map(D => n_346, E => n_889, Q => FE_OFN117_snake_output22_4);
  S_S_reg_22_5 : LHQD1BWP7T port map(D => n_347, E => n_889, Q => FE_OFN151_snake_output22_5);
  S_S_reg_23_0 : LHQD1BWP7T port map(D => n_369, E => n_888, Q => FE_OFN133_snake_output23_0);
  S_S_reg_23_1 : LHQD1BWP7T port map(D => n_368, E => n_888, Q => FE_OFN131_snake_output23_1);
  S_S_reg_23_2 : LHQD1BWP7T port map(D => n_366, E => n_888, Q => FE_OFN128_snake_output23_2);
  S_S_reg_23_3 : LHQD1BWP7T port map(D => n_341, E => n_888, Q => FE_OFN132_snake_output23_3);
  S_S_reg_23_4 : LHQD1BWP7T port map(D => n_365, E => n_888, Q => FE_OFN130_snake_output23_4);
  S_S_reg_23_5 : LHQD1BWP7T port map(D => n_364, E => n_888, Q => n_1053);
  S_S_reg_24_0 : LHQD1BWP7T port map(D => n_362, E => n_890, Q => FE_OFN155_snake_output24_0);
  S_S_reg_24_1 : LHQD1BWP7T port map(D => n_361, E => n_890, Q => FE_OFN158_snake_output24_1);
  S_S_reg_24_2 : LHQD1BWP7T port map(D => n_351, E => n_890, Q => FE_OFN157_snake_output24_2);
  S_S_reg_24_3 : LHQD1BWP7T port map(D => n_358, E => n_890, Q => FE_OFN154_snake_output24_3);
  S_S_reg_24_4 : LHQD1BWP7T port map(D => n_359, E => n_890, Q => FE_OFN156_snake_output24_4);
  S_S_reg_24_5 : LHQD1BWP7T port map(D => n_357, E => n_890, Q => FE_OFN159_snake_output24_5);
  corner_check_reg_5 : LNQD1BWP7T port map(D => n_1037, EN => n_530, Q => corner_check(5));
  corner_count_reg_0 : LNQD1BWP7T port map(D => n_451, EN => n_470, Q => corner_count(0));
  corner_count_reg_1 : LNQD1BWP7T port map(D => n_251, EN => n_470, Q => corner_count(1));
  corner_count_reg_2 : LNQD1BWP7T port map(D => n_269, EN => n_470, Q => corner_count(2));
  corner_count_reg_3 : LNQD1BWP7T port map(D => n_268, EN => n_470, Q => corner_count(3));
  corner_count_reg_4 : LNQD1BWP7T port map(D => n_270, EN => n_470, Q => corner_count(4));
  corner_count_reg_5 : LNQD1BWP7T port map(D => n_267, EN => n_470, Q => corner_count(5));
  corner_count_reg_6 : LNQD1BWP7T port map(D => n_266, EN => n_470, Q => corner_count(6));
  corner_count_reg_7 : LNQD1BWP7T port map(D => n_265, EN => n_470, Q => corner_count(7));
  corner_count_reg_8 : LNQD1BWP7T port map(D => n_264, EN => n_470, Q => corner_count(8));
  corner_count_reg_9 : LNQD1BWP7T port map(D => n_272, EN => n_470, Q => corner_count(9));
  corner_count_reg_10 : LNQD1BWP7T port map(D => n_271, EN => n_470, Q => corner_count(10));
  corner_count_reg_11 : LNQD1BWP7T port map(D => n_262, EN => n_470, Q => corner_count(11));
  corner_count_reg_12 : LNQD1BWP7T port map(D => n_250, EN => n_470, Q => corner_count(12));
  corner_count_reg_13 : LNQD1BWP7T port map(D => n_261, EN => n_470, Q => corner_count(13));
  corner_count_reg_14 : LNQD1BWP7T port map(D => n_247, EN => n_470, Q => corner_count(14));
  corner_count_reg_15 : LNQD1BWP7T port map(D => n_242, EN => n_470, Q => corner_count(15));
  corner_count_reg_16 : LNQD1BWP7T port map(D => n_241, EN => n_470, Q => corner_count(16));
  corner_count_reg_17 : LNQD1BWP7T port map(D => n_253, EN => n_470, Q => corner_count(17));
  corner_count_reg_18 : LNQD1BWP7T port map(D => n_260, EN => n_470, Q => corner_count(18));
  corner_count_reg_19 : LNQD1BWP7T port map(D => n_259, EN => n_470, Q => corner_count(19));
  corner_count_reg_20 : LNQD1BWP7T port map(D => n_244, EN => n_470, Q => corner_count(20));
  corner_count_reg_21 : LNQD1BWP7T port map(D => n_248, EN => n_470, Q => corner_count(21));
  corner_count_reg_22 : LNQD1BWP7T port map(D => n_263, EN => n_470, Q => corner_count(22));
  corner_count_reg_23 : LNQD1BWP7T port map(D => n_258, EN => n_470, Q => corner_count(23));
  corner_count_reg_24 : LNQD1BWP7T port map(D => n_243, EN => n_470, Q => corner_count(24));
  corner_count_reg_25 : LNQD1BWP7T port map(D => n_245, EN => n_470, Q => corner_count(25));
  corner_count_reg_26 : LNQD1BWP7T port map(D => n_257, EN => n_470, Q => corner_count(26));
  corner_count_reg_27 : LNQD1BWP7T port map(D => n_256, EN => n_470, Q => corner_count(27));
  corner_count_reg_28 : LNQD1BWP7T port map(D => n_246, EN => n_470, Q => corner_count(28));
  corner_count_reg_29 : LNQD1BWP7T port map(D => n_249, EN => n_470, Q => corner_count(29));
  corner_count_reg_30 : LNQD1BWP7T port map(D => n_255, EN => n_470, Q => corner_count(30));
  corner_count_reg_31 : LNQD1BWP7T port map(D => n_252, EN => n_470, Q => corner_count(31));
  new_N_reg_1 : LNQD1BWP7T port map(D => n_1617, EN => FE_OFN2_n_1651, Q => new_N(1));
  new_N_reg_2 : LNQD1BWP7T port map(D => n_1616, EN => FE_OFN2_n_1651, Q => new_N(2));
  new_N_reg_3 : LNQD1BWP7T port map(D => n_1615, EN => FE_OFN2_n_1651, Q => new_N(3));
  new_N_reg_4 : LNQD1BWP7T port map(D => n_1614, EN => FE_OFN2_n_1651, Q => new_N(4));
  new_N_reg_5 : LNQD1BWP7T port map(D => n_1613, EN => FE_OFN2_n_1651, Q => new_N(5));
  new_N_reg_6 : LNQD1BWP7T port map(D => n_1612, EN => FE_OFN2_n_1651, Q => new_N(6));
  new_N_reg_7 : LNQD1BWP7T port map(D => n_1611, EN => FE_OFN2_n_1651, Q => new_N(7));
  new_N_reg_8 : LNQD1BWP7T port map(D => n_1610, EN => FE_OFN2_n_1651, Q => new_N(8));
  new_N_reg_9 : LNQD1BWP7T port map(D => n_1609, EN => FE_OFN2_n_1651, Q => new_N(9));
  new_N_reg_10 : LNQD1BWP7T port map(D => n_1608, EN => FE_OFN2_n_1651, Q => new_N(10));
  new_N_reg_11 : LNQD1BWP7T port map(D => n_1607, EN => FE_OFN2_n_1651, Q => new_N(11));
  new_N_reg_12 : LNQD1BWP7T port map(D => n_1606, EN => FE_OFN2_n_1651, Q => new_N(12));
  new_N_reg_13 : LNQD1BWP7T port map(D => n_1605, EN => FE_OFN2_n_1651, Q => new_N(13));
  new_N_reg_14 : LNQD1BWP7T port map(D => n_1604, EN => FE_OFN2_n_1651, Q => new_N(14));
  new_N_reg_15 : LNQD1BWP7T port map(D => n_1603, EN => FE_OFN2_n_1651, Q => new_N(15));
  new_N_reg_16 : LNQD1BWP7T port map(D => n_1602, EN => FE_OFN2_n_1651, Q => new_N(16));
  new_N_reg_17 : LNQD1BWP7T port map(D => n_1601, EN => FE_OFN2_n_1651, Q => new_N(17));
  new_N_reg_18 : LNQD1BWP7T port map(D => n_1600, EN => FE_OFN2_n_1651, Q => new_N(18));
  new_N_reg_19 : LNQD1BWP7T port map(D => n_1599, EN => FE_OFN2_n_1651, Q => new_N(19));
  new_N_reg_20 : LNQD1BWP7T port map(D => n_1598, EN => FE_OFN2_n_1651, Q => new_N(20));
  new_N_reg_21 : LNQD1BWP7T port map(D => n_1597, EN => FE_OFN2_n_1651, Q => new_N(21));
  new_N_reg_22 : LNQD1BWP7T port map(D => n_1596, EN => FE_OFN2_n_1651, Q => new_N(22));
  new_N_reg_23 : LNQD1BWP7T port map(D => n_1595, EN => FE_OFN2_n_1651, Q => new_N(23));
  new_N_reg_24 : LNQD1BWP7T port map(D => n_1594, EN => FE_OFN2_n_1651, Q => new_N(24));
  new_N_reg_25 : LNQD1BWP7T port map(D => n_1593, EN => FE_OFN2_n_1651, Q => new_N(25));
  new_N_reg_26 : LNQD1BWP7T port map(D => n_1592, EN => FE_OFN2_n_1651, Q => new_N(26));
  new_N_reg_27 : LNQD1BWP7T port map(D => n_1591, EN => FE_OFN2_n_1651, Q => new_N(27));
  new_N_reg_28 : LNQD1BWP7T port map(D => n_1590, EN => FE_OFN2_n_1651, Q => new_N(28));
  new_N_reg_29 : LNQD1BWP7T port map(D => n_1589, EN => FE_OFN2_n_1651, Q => new_N(29));
  new_N_reg_30 : LNQD1BWP7T port map(D => n_1588, EN => FE_OFN2_n_1651, Q => new_N(30));
  new_N_reg_31 : LNQD1BWP7T port map(D => n_1587, EN => FE_OFN2_n_1651, Q => new_N(31));
  new_corner_count_reg_1 : LHQD1BWP7T port map(D => n_1648, E => FE_OFN0_n_1657, Q => new_corner_count(1));
  new_corner_count_reg_2 : LHQD1BWP7T port map(D => n_1647, E => FE_OFN0_n_1657, Q => new_corner_count(2));
  new_corner_count_reg_3 : LHQD1BWP7T port map(D => n_1646, E => FE_OFN0_n_1657, Q => new_corner_count(3));
  new_corner_count_reg_4 : LHQD1BWP7T port map(D => n_1645, E => FE_OFN0_n_1657, Q => new_corner_count(4));
  new_corner_count_reg_5 : LHQD1BWP7T port map(D => n_1644, E => FE_OFN0_n_1657, Q => new_corner_count(5));
  new_corner_count_reg_6 : LHQD1BWP7T port map(D => n_1643, E => FE_OFN0_n_1657, Q => new_corner_count(6));
  new_corner_count_reg_7 : LHQD1BWP7T port map(D => n_1642, E => FE_OFN0_n_1657, Q => new_corner_count(7));
  new_corner_count_reg_8 : LHQD1BWP7T port map(D => n_1641, E => FE_OFN0_n_1657, Q => new_corner_count(8));
  new_corner_count_reg_9 : LHQD1BWP7T port map(D => n_1640, E => FE_OFN0_n_1657, Q => new_corner_count(9));
  new_corner_count_reg_10 : LHQD1BWP7T port map(D => n_1639, E => FE_OFN0_n_1657, Q => new_corner_count(10));
  new_corner_count_reg_11 : LHQD1BWP7T port map(D => n_1638, E => FE_OFN0_n_1657, Q => new_corner_count(11));
  new_corner_count_reg_12 : LHQD1BWP7T port map(D => n_1637, E => FE_OFN0_n_1657, Q => new_corner_count(12));
  new_corner_count_reg_13 : LHQD1BWP7T port map(D => n_1636, E => FE_OFN0_n_1657, Q => new_corner_count(13));
  new_corner_count_reg_14 : LHQD1BWP7T port map(D => n_1635, E => FE_OFN0_n_1657, Q => new_corner_count(14));
  new_corner_count_reg_15 : LHQD1BWP7T port map(D => n_1634, E => FE_OFN0_n_1657, Q => new_corner_count(15));
  new_corner_count_reg_16 : LHQD1BWP7T port map(D => n_1633, E => FE_OFN0_n_1657, Q => new_corner_count(16));
  new_corner_count_reg_17 : LHQD1BWP7T port map(D => n_1632, E => FE_OFN0_n_1657, Q => new_corner_count(17));
  new_corner_count_reg_18 : LHQD1BWP7T port map(D => n_1631, E => FE_OFN0_n_1657, Q => new_corner_count(18));
  new_corner_count_reg_19 : LHQD1BWP7T port map(D => n_1630, E => FE_OFN0_n_1657, Q => new_corner_count(19));
  new_corner_count_reg_20 : LHQD1BWP7T port map(D => n_1629, E => FE_OFN0_n_1657, Q => new_corner_count(20));
  new_corner_count_reg_21 : LHQD1BWP7T port map(D => n_1628, E => FE_OFN0_n_1657, Q => new_corner_count(21));
  new_corner_count_reg_22 : LHQD1BWP7T port map(D => n_1627, E => FE_OFN0_n_1657, Q => new_corner_count(22));
  new_corner_count_reg_23 : LHQD1BWP7T port map(D => n_1626, E => n_1657, Q => new_corner_count(23));
  new_corner_count_reg_24 : LHQD1BWP7T port map(D => n_1625, E => n_1657, Q => new_corner_count(24));
  new_corner_count_reg_25 : LHQD1BWP7T port map(D => n_1624, E => n_1657, Q => new_corner_count(25));
  new_corner_count_reg_26 : LHQD1BWP7T port map(D => n_1623, E => n_1657, Q => new_corner_count(26));
  new_corner_count_reg_27 : LHQD1BWP7T port map(D => n_1622, E => n_1657, Q => new_corner_count(27));
  new_corner_count_reg_28 : LHQD1BWP7T port map(D => n_1621, E => n_1657, Q => new_corner_count(28));
  new_corner_count_reg_29 : LHQD1BWP7T port map(D => n_1620, E => n_1657, Q => new_corner_count(29));
  new_corner_count_reg_30 : LHQD1BWP7T port map(D => n_1619, E => n_1657, Q => new_corner_count(30));
  new_corner_count_reg_31 : LHQD1BWP7T port map(D => n_1618, E => n_1657, Q => new_corner_count(31));
  new_state_reg_0 : LHQD1BWP7T port map(D => n_1040, E => n_1649, Q => new_state(0));
  new_state_reg_1 : LHQD1BWP7T port map(D => n_1041, E => n_1649, Q => new_state(1));
  shift0_reg_0 : LHQD1BWP7T port map(D => snake_output0(0), E => n_1657, Q => shift0(0));
  shift0_reg_1 : LHQD1BWP7T port map(D => snake_output0(1), E => n_1657, Q => shift0(1));
  shift0_reg_2 : LHQD1BWP7T port map(D => snake_output0(2), E => n_1657, Q => shift0(2));
  shift0_reg_3 : LHQD1BWP7T port map(D => snake_output0(3), E => n_1657, Q => shift0(3));
  shift0_reg_4 : LHQD1BWP7T port map(D => snake_output0(4), E => n_1657, Q => shift0(4));
  shift0_reg_5 : LHQD1BWP7T port map(D => snake_output0(5), E => n_1657, Q => shift0(5));
  shift1_reg_0 : LHQD1BWP7T port map(D => snake_output1(0), E => n_1657, Q => shift1(0));
  shift1_reg_1 : LHQD1BWP7T port map(D => snake_output1(1), E => n_1657, Q => shift1(1));
  shift1_reg_2 : LHQD1BWP7T port map(D => snake_output1(2), E => n_1657, Q => shift1(2));
  shift1_reg_3 : LHQD1BWP7T port map(D => snake_output1(3), E => n_1657, Q => shift1(3));
  shift1_reg_4 : LHQD1BWP7T port map(D => snake_output1(4), E => n_1657, Q => shift1(4));
  shift1_reg_5 : LHQD1BWP7T port map(D => snake_output1(5), E => n_1657, Q => shift1(5));
  shift2_reg_0 : LHQD1BWP7T port map(D => snake_output2(0), E => FE_OFN0_n_1657, Q => shift2(0));
  shift2_reg_1 : LHQD1BWP7T port map(D => snake_output2(1), E => n_1657, Q => shift2(1));
  shift2_reg_2 : LHQD1BWP7T port map(D => snake_output2(2), E => FE_OFN0_n_1657, Q => shift2(2));
  shift2_reg_3 : LHQD1BWP7T port map(D => snake_output2(3), E => n_1657, Q => shift2(3));
  shift2_reg_4 : LHQD1BWP7T port map(D => snake_output2(4), E => n_1657, Q => shift2(4));
  shift2_reg_5 : LHQD1BWP7T port map(D => snake_output2(5), E => FE_OFN0_n_1657, Q => shift2(5));
  shift3_reg_0 : LHQD1BWP7T port map(D => snake_output3(0), E => FE_OFN0_n_1657, Q => shift3(0));
  shift3_reg_1 : LHQD1BWP7T port map(D => snake_output3(1), E => n_1657, Q => shift3(1));
  shift3_reg_2 : LHQD1BWP7T port map(D => snake_output3(2), E => n_1657, Q => shift3(2));
  shift3_reg_3 : LHQD1BWP7T port map(D => snake_output3(3), E => n_1657, Q => shift3(3));
  shift3_reg_4 : LHQD1BWP7T port map(D => snake_output3(4), E => n_1657, Q => shift3(4));
  shift3_reg_5 : LHQD1BWP7T port map(D => snake_output3(5), E => FE_OFN0_n_1657, Q => shift3(5));
  shift4_reg_0 : LHQD1BWP7T port map(D => snake_output4(0), E => FE_OFN0_n_1657, Q => shift4(0));
  shift4_reg_1 : LHQD1BWP7T port map(D => snake_output4(1), E => FE_OFN0_n_1657, Q => shift4(1));
  shift4_reg_2 : LHQD1BWP7T port map(D => snake_output4(2), E => FE_OFN0_n_1657, Q => shift4(2));
  shift4_reg_3 : LHQD1BWP7T port map(D => snake_output4(3), E => n_1657, Q => shift4(3));
  shift4_reg_4 : LHQD1BWP7T port map(D => snake_output4(4), E => FE_OFN0_n_1657, Q => shift4(4));
  shift4_reg_5 : LHQD1BWP7T port map(D => n_1167, E => FE_OFN0_n_1657, Q => shift4(5));
  shift5_reg_0 : LHQD1BWP7T port map(D => snake_output5(0), E => FE_OFN0_n_1657, Q => shift5(0));
  shift5_reg_1 : LHQD1BWP7T port map(D => snake_output5(1), E => FE_OFN0_n_1657, Q => shift5(1));
  shift5_reg_2 : LHQD1BWP7T port map(D => snake_output5(2), E => FE_OFN0_n_1657, Q => shift5(2));
  shift5_reg_3 : LHQD1BWP7T port map(D => snake_output5(3), E => FE_OFN0_n_1657, Q => shift5(3));
  shift5_reg_4 : LHQD1BWP7T port map(D => snake_output5(4), E => FE_OFN0_n_1657, Q => shift5(4));
  shift5_reg_5 : LHQD1BWP7T port map(D => snake_output5(5), E => FE_OFN0_n_1657, Q => shift5(5));
  shift6_reg_0 : LHQD1BWP7T port map(D => snake_output6(0), E => FE_OFN0_n_1657, Q => shift6(0));
  shift6_reg_1 : LHQD1BWP7T port map(D => snake_output6(1), E => FE_OFN0_n_1657, Q => shift6(1));
  shift6_reg_2 : LHQD1BWP7T port map(D => snake_output6(2), E => FE_OFN0_n_1657, Q => shift6(2));
  shift6_reg_3 : LHQD1BWP7T port map(D => snake_output6(3), E => FE_OFN0_n_1657, Q => shift6(3));
  shift6_reg_4 : LHQD1BWP7T port map(D => snake_output6(4), E => FE_OFN0_n_1657, Q => shift6(4));
  shift6_reg_5 : LHQD1BWP7T port map(D => snake_output6(5), E => FE_OFN0_n_1657, Q => shift6(5));
  shift7_reg_0 : LHQD1BWP7T port map(D => snake_output7(0), E => FE_OFN0_n_1657, Q => shift7(0));
  shift7_reg_1 : LHQD1BWP7T port map(D => snake_output7(1), E => FE_OFN0_n_1657, Q => shift7(1));
  shift7_reg_2 : LHQD1BWP7T port map(D => snake_output7(2), E => FE_OFN0_n_1657, Q => shift7(2));
  shift7_reg_3 : LHQD1BWP7T port map(D => snake_output7(3), E => FE_OFN0_n_1657, Q => shift7(3));
  shift7_reg_4 : LHQD1BWP7T port map(D => snake_output7(4), E => FE_OFN0_n_1657, Q => shift7(4));
  shift7_reg_5 : LHQD1BWP7T port map(D => snake_output7(5), E => FE_OFN0_n_1657, Q => shift7(5));
  shift8_reg_0 : LHQD1BWP7T port map(D => snake_output8(0), E => FE_OFN0_n_1657, Q => shift8(0));
  shift8_reg_1 : LHQD1BWP7T port map(D => snake_output8(1), E => FE_OFN0_n_1657, Q => shift8(1));
  shift8_reg_2 : LHQD1BWP7T port map(D => snake_output8(2), E => FE_OFN0_n_1657, Q => shift8(2));
  shift8_reg_3 : LHQD1BWP7T port map(D => snake_output8(3), E => FE_OFN0_n_1657, Q => shift8(3));
  shift8_reg_4 : LHQD1BWP7T port map(D => snake_output8(4), E => FE_OFN0_n_1657, Q => shift8(4));
  shift8_reg_5 : LHQD1BWP7T port map(D => snake_output8(5), E => FE_OFN0_n_1657, Q => shift8(5));
  shift9_reg_0 : LHQD1BWP7T port map(D => snake_output9(0), E => FE_OFN0_n_1657, Q => shift9(0));
  shift9_reg_1 : LHQD1BWP7T port map(D => snake_output9(1), E => FE_OFN1_n_1657, Q => shift9(1));
  shift9_reg_2 : LHQD1BWP7T port map(D => snake_output9(2), E => FE_OFN1_n_1657, Q => shift9(2));
  shift9_reg_3 : LHQD1BWP7T port map(D => snake_output9(3), E => FE_OFN1_n_1657, Q => shift9(3));
  shift9_reg_4 : LHQD1BWP7T port map(D => snake_output9(4), E => FE_OFN1_n_1657, Q => shift9(4));
  shift9_reg_5 : LHQD1BWP7T port map(D => snake_output9(5), E => FE_OFN0_n_1657, Q => shift9(5));
  shift10_reg_0 : LHQD1BWP7T port map(D => snake_output10(0), E => FE_OFN1_n_1657, Q => shift10(0));
  shift10_reg_1 : LHQD1BWP7T port map(D => snake_output10(1), E => FE_OFN1_n_1657, Q => shift10(1));
  shift10_reg_2 : LHQD1BWP7T port map(D => snake_output10(2), E => FE_OFN1_n_1657, Q => shift10(2));
  shift10_reg_3 : LHQD1BWP7T port map(D => snake_output10(3), E => FE_OFN1_n_1657, Q => shift10(3));
  shift10_reg_4 : LHQD1BWP7T port map(D => snake_output10(4), E => FE_OFN1_n_1657, Q => shift10(4));
  shift10_reg_5 : LHQD1BWP7T port map(D => snake_output10(5), E => FE_OFN0_n_1657, Q => shift10(5));
  shift11_reg_0 : LHQD1BWP7T port map(D => snake_output11(0), E => FE_OFN1_n_1657, Q => shift11(0));
  shift11_reg_1 : LHQD1BWP7T port map(D => snake_output11(1), E => FE_OFN1_n_1657, Q => shift11(1));
  shift11_reg_2 : LHQD1BWP7T port map(D => snake_output11(2), E => FE_OFN1_n_1657, Q => shift11(2));
  shift11_reg_3 : LHQD1BWP7T port map(D => snake_output11(3), E => FE_OFN1_n_1657, Q => shift11(3));
  shift11_reg_4 : LHQD1BWP7T port map(D => snake_output11(4), E => FE_OFN1_n_1657, Q => shift11(4));
  shift11_reg_5 : LHQD1BWP7T port map(D => snake_output11(5), E => FE_OFN0_n_1657, Q => shift11(5));
  shift12_reg_0 : LHQD1BWP7T port map(D => snake_output12(0), E => FE_OFN1_n_1657, Q => shift12(0));
  shift12_reg_1 : LHQD1BWP7T port map(D => snake_output12(1), E => FE_OFN1_n_1657, Q => shift12(1));
  shift12_reg_2 : LHQD1BWP7T port map(D => snake_output12(2), E => FE_OFN1_n_1657, Q => shift12(2));
  shift12_reg_3 : LHQD1BWP7T port map(D => snake_output12(3), E => FE_OFN1_n_1657, Q => shift12(3));
  shift12_reg_4 : LHQD1BWP7T port map(D => snake_output12(4), E => FE_OFN1_n_1657, Q => shift12(4));
  shift12_reg_5 : LHQD1BWP7T port map(D => snake_output12(5), E => FE_OFN0_n_1657, Q => shift12(5));
  shift13_reg_0 : LHQD1BWP7T port map(D => snake_output13(0), E => FE_OFN1_n_1657, Q => shift13(0));
  shift13_reg_1 : LHQD1BWP7T port map(D => snake_output13(1), E => FE_OFN1_n_1657, Q => shift13(1));
  shift13_reg_2 : LHQD1BWP7T port map(D => snake_output13(2), E => FE_OFN1_n_1657, Q => shift13(2));
  shift13_reg_3 : LHQD1BWP7T port map(D => snake_output13(3), E => FE_OFN1_n_1657, Q => shift13(3));
  shift13_reg_4 : LHQD1BWP7T port map(D => snake_output13(4), E => FE_OFN1_n_1657, Q => shift13(4));
  shift13_reg_5 : LHQD1BWP7T port map(D => snake_output13(5), E => FE_OFN0_n_1657, Q => shift13(5));
  shift14_reg_0 : LHQD1BWP7T port map(D => snake_output14(0), E => FE_OFN0_n_1657, Q => shift14(0));
  shift14_reg_1 : LHQD1BWP7T port map(D => snake_output14(1), E => FE_OFN1_n_1657, Q => shift14(1));
  shift14_reg_2 : LHQD1BWP7T port map(D => snake_output14(2), E => FE_OFN1_n_1657, Q => shift14(2));
  shift14_reg_3 : LHQD1BWP7T port map(D => snake_output14(3), E => FE_OFN1_n_1657, Q => shift14(3));
  shift14_reg_4 : LHQD1BWP7T port map(D => snake_output14(4), E => FE_OFN1_n_1657, Q => shift14(4));
  shift14_reg_5 : LHQD1BWP7T port map(D => snake_output14(5), E => FE_OFN0_n_1657, Q => shift14(5));
  shift15_reg_0 : LHQD1BWP7T port map(D => snake_output15(0), E => FE_OFN1_n_1657, Q => shift15(0));
  shift15_reg_1 : LHQD1BWP7T port map(D => snake_output15(1), E => FE_OFN1_n_1657, Q => shift15(1));
  shift15_reg_2 : LHQD1BWP7T port map(D => snake_output15(2), E => FE_OFN1_n_1657, Q => shift15(2));
  shift15_reg_3 : LHQD1BWP7T port map(D => snake_output15(3), E => FE_OFN1_n_1657, Q => shift15(3));
  shift15_reg_4 : LHQD1BWP7T port map(D => snake_output15(4), E => FE_OFN1_n_1657, Q => shift15(4));
  shift15_reg_5 : LHQD1BWP7T port map(D => snake_output15(5), E => FE_OFN0_n_1657, Q => shift15(5));
  shift16_reg_0 : LHQD1BWP7T port map(D => snake_output16(0), E => FE_OFN1_n_1657, Q => shift16(0));
  shift16_reg_1 : LHQD1BWP7T port map(D => snake_output16(1), E => FE_OFN1_n_1657, Q => shift16(1));
  shift16_reg_2 : LHQD1BWP7T port map(D => snake_output16(2), E => FE_OFN1_n_1657, Q => shift16(2));
  shift16_reg_3 : LHQD1BWP7T port map(D => snake_output16(3), E => FE_OFN1_n_1657, Q => shift16(3));
  shift16_reg_4 : LHQD1BWP7T port map(D => snake_output16(4), E => FE_OFN1_n_1657, Q => shift16(4));
  shift16_reg_5 : LHQD1BWP7T port map(D => snake_output16(5), E => FE_OFN0_n_1657, Q => shift16(5));
  shift17_reg_0 : LHQD1BWP7T port map(D => snake_output17(0), E => FE_OFN1_n_1657, Q => shift17(0));
  shift17_reg_1 : LHQD1BWP7T port map(D => snake_output17(1), E => FE_OFN1_n_1657, Q => shift17(1));
  shift17_reg_2 : LHQD1BWP7T port map(D => snake_output17(2), E => FE_OFN1_n_1657, Q => shift17(2));
  shift17_reg_3 : LHQD1BWP7T port map(D => snake_output17(3), E => FE_OFN1_n_1657, Q => shift17(3));
  shift17_reg_4 : LHQD1BWP7T port map(D => snake_output17(4), E => FE_OFN1_n_1657, Q => shift17(4));
  shift17_reg_5 : LHQD1BWP7T port map(D => snake_output17(5), E => FE_OFN0_n_1657, Q => shift17(5));
  shift18_reg_0 : LHQD1BWP7T port map(D => snake_output18(0), E => FE_OFN1_n_1657, Q => shift18(0));
  shift18_reg_1 : LHQD1BWP7T port map(D => snake_output18(1), E => FE_OFN1_n_1657, Q => shift18(1));
  shift18_reg_2 : LHQD1BWP7T port map(D => snake_output18(2), E => FE_OFN1_n_1657, Q => shift18(2));
  shift18_reg_3 : LHQD1BWP7T port map(D => snake_output18(3), E => FE_OFN1_n_1657, Q => shift18(3));
  shift18_reg_4 : LHQD1BWP7T port map(D => snake_output18(4), E => FE_OFN1_n_1657, Q => shift18(4));
  shift18_reg_5 : LHQD1BWP7T port map(D => snake_output18(5), E => FE_OFN0_n_1657, Q => shift18(5));
  shift19_reg_0 : LHQD1BWP7T port map(D => snake_output19(0), E => FE_OFN1_n_1657, Q => shift19(0));
  shift19_reg_1 : LHQD1BWP7T port map(D => snake_output19(1), E => FE_OFN1_n_1657, Q => shift19(1));
  shift19_reg_2 : LHQD1BWP7T port map(D => snake_output19(2), E => FE_OFN1_n_1657, Q => shift19(2));
  shift19_reg_3 : LHQD1BWP7T port map(D => snake_output19(3), E => FE_OFN1_n_1657, Q => shift19(3));
  shift19_reg_4 : LHQD1BWP7T port map(D => snake_output19(4), E => FE_OFN1_n_1657, Q => shift19(4));
  shift19_reg_5 : LHQD1BWP7T port map(D => snake_output19(5), E => FE_OFN0_n_1657, Q => shift19(5));
  shift20_reg_0 : LHQD1BWP7T port map(D => snake_output20(0), E => FE_OFN1_n_1657, Q => shift20(0));
  shift20_reg_1 : LHQD1BWP7T port map(D => snake_output20(1), E => FE_OFN1_n_1657, Q => shift20(1));
  shift20_reg_2 : LHQD1BWP7T port map(D => snake_output20(2), E => FE_OFN1_n_1657, Q => shift20(2));
  shift20_reg_3 : LHQD1BWP7T port map(D => snake_output20(3), E => FE_OFN1_n_1657, Q => shift20(3));
  shift20_reg_4 : LHQD1BWP7T port map(D => snake_output20(4), E => FE_OFN1_n_1657, Q => shift20(4));
  shift20_reg_5 : LHQD1BWP7T port map(D => snake_output20(5), E => FE_OFN0_n_1657, Q => shift20(5));
  shift21_reg_0 : LHQD1BWP7T port map(D => snake_output21(0), E => FE_OFN1_n_1657, Q => shift21(0));
  shift21_reg_1 : LHQD1BWP7T port map(D => snake_output21(1), E => FE_OFN1_n_1657, Q => shift21(1));
  shift21_reg_2 : LHQD1BWP7T port map(D => snake_output21(2), E => FE_OFN1_n_1657, Q => shift21(2));
  shift21_reg_3 : LHQD1BWP7T port map(D => snake_output21(3), E => FE_OFN1_n_1657, Q => shift21(3));
  shift21_reg_4 : LHQD1BWP7T port map(D => snake_output21(4), E => FE_OFN1_n_1657, Q => shift21(4));
  shift21_reg_5 : LHQD1BWP7T port map(D => snake_output21(5), E => FE_OFN0_n_1657, Q => shift21(5));
  shift22_reg_0 : LHQD1BWP7T port map(D => snake_output22(0), E => FE_OFN1_n_1657, Q => shift22(0));
  shift22_reg_1 : LHQD1BWP7T port map(D => snake_output22(1), E => FE_OFN1_n_1657, Q => shift22(1));
  shift22_reg_2 : LHQD1BWP7T port map(D => snake_output22(2), E => FE_OFN1_n_1657, Q => shift22(2));
  shift22_reg_3 : LHQD1BWP7T port map(D => snake_output22(3), E => FE_OFN1_n_1657, Q => shift22(3));
  shift22_reg_4 : LHQD1BWP7T port map(D => snake_output22(4), E => FE_OFN1_n_1657, Q => shift22(4));
  shift22_reg_5 : LHQD1BWP7T port map(D => snake_output22(5), E => FE_OFN0_n_1657, Q => shift22(5));
  shift23_reg_0 : LHQD1BWP7T port map(D => snake_output23(0), E => FE_OFN1_n_1657, Q => shift23(0));
  shift23_reg_1 : LHQD1BWP7T port map(D => snake_output23(1), E => FE_OFN1_n_1657, Q => shift23(1));
  shift23_reg_2 : LHQD1BWP7T port map(D => snake_output23(2), E => FE_OFN1_n_1657, Q => shift23(2));
  shift23_reg_3 : LHQD1BWP7T port map(D => snake_output23(3), E => FE_OFN1_n_1657, Q => shift23(3));
  shift23_reg_4 : LHQD1BWP7T port map(D => snake_output23(4), E => FE_OFN1_n_1657, Q => shift23(4));
  shift23_reg_5 : LHQD1BWP7T port map(D => n_1053, E => FE_OFN0_n_1657, Q => shift23(5));
  snake_list_reg_1 : LHQD1BWP7T port map(D => n_992, E => n_1652, Q => FE_OFN175_snake_list_1);
  snake_list_reg_2 : LHQD1BWP7T port map(D => n_991, E => n_1652, Q => FE_OFN168_snake_list_2);
  snake_list_reg_3 : LHQD1BWP7T port map(D => n_990, E => n_1652, Q => FE_OFN173_snake_list_3);
  snake_list_reg_4 : LHQD1BWP7T port map(D => n_989, E => n_1652, Q => FE_OFN167_snake_list_4);
  snake_list_reg_5 : LHQD1BWP7T port map(D => n_988, E => n_1652, Q => FE_OFN171_snake_list_5);
  snake_list_reg_6 : LHQD1BWP7T port map(D => n_952, E => n_1652, Q => FE_OFN160_snake_list_6);
  snake_list_reg_7 : LHQD1BWP7T port map(D => n_1018, E => n_1652, Q => FE_OFN164_snake_list_7);
  snake_list_reg_8 : LHQD1BWP7T port map(D => n_1030, E => n_1652, Q => FE_OFN169_snake_list_8);
  snake_list_reg_9 : LHQD1BWP7T port map(D => n_1017, E => n_1652, Q => FE_OFN162_snake_list_9);
  snake_list_reg_10 : LHQD1BWP7T port map(D => n_1023, E => n_1652, Q => FE_OFN172_snake_list_10);
  snake_list_reg_11 : LHQD1BWP7T port map(D => n_1029, E => n_1652, Q => FE_OFN165_snake_list_11);
  snake_list_reg_12 : LHQD1BWP7T port map(D => n_1028, E => n_1652, Q => FE_OFN163_snake_list_12);
  snake_list_reg_13 : LHQD1BWP7T port map(D => n_1026, E => n_1652, Q => FE_OFN174_snake_list_13);
  snake_list_reg_14 : LHQD1BWP7T port map(D => n_1016, E => n_1652, Q => FE_OFN161_snake_list_14);
  snake_list_reg_15 : LHQD1BWP7T port map(D => n_1031, E => n_1652, Q => FE_OFN170_snake_list_15);
  snake_list_reg_16 : LHQD1BWP7T port map(D => n_1025, E => n_1652, Q => FE_OFN166_snake_list_16);
  state_reg_1 : DFKCNQD1BWP7T port map(CN => new_state(1), CP => CTS_6, D => n_157, Q => state(1));
  state_reg_3 : DFKCNQD1BWP7T port map(CN => new_state(3), CP => CTS_6, D => n_157, Q => state(3));
  state_reg_4 : DFKCNQD1BWP7T port map(CN => new_state(4), CP => CTS_6, D => n_157, Q => state(4));
  g29160 : OR4D0BWP7T port map(A1 => n_1736, A2 => n_1748, A3 => n_236, A4 => n_1039, Z => n_1041);
  g29161 : NR4D0BWP7T port map(A1 => n_1039, A2 => n_236, A3 => n_676, A4 => n_1657, ZN => n_1040);
  g29162 : NR3D0BWP7T port map(A1 => n_1032, A2 => n_1038, A3 => n_1022, ZN => n_1039);
  g29164 : AO211D0BWP7T port map(A1 => n_1036, A2 => n_419, B => n_1035, C => n_1021, Z => n_1038);
  g29165 : OAI211D0BWP7T port map(A1 => n_221, A2 => n_472, B => n_1034, C => n_494, ZN => n_1037);
  g29166 : INR4D0BWP7T port map(A1 => n_1024, B1 => corner_count(11), B2 => corner_count(12), B3 => corner_count(4), ZN => n_1036);
  g29167 : OAI221D0BWP7T port map(A1 => n_1012, A2 => new_tail(2), B1 => new_tail(0), B2 => n_1013, C => n_1033, ZN => n_1035);
  g29168 : OA221D0BWP7T port map(A1 => n_473, A2 => n_213, B1 => n_440, B2 => n_471, C => n_1027, Z => n_1034);
  g29176 : AOI221D0BWP7T port map(A1 => n_1012, A2 => new_tail(2), B1 => n_1013, B2 => new_tail(0), C => n_1020, ZN => n_1033);
  g29177 : OAI211D0BWP7T port map(A1 => new_tail(4), A2 => n_1015, B => n_1571, C => n_1019, ZN => n_1032);
  g29178 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_984, B => n_1003, C => n_456, ZN => n_1031);
  g29181 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_995, B => n_1007, C => n_444, ZN => n_1030);
  g29182 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_987, B => n_1002, C => n_450, ZN => n_1029);
  g29183 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_976, B => n_1001, C => n_454, ZN => n_1028);
  g29185 : AN4D1BWP7T port map(A1 => n_1000, A2 => n_679, A3 => n_526, A4 => n_490, Z => n_1027);
  g29186 : OAI211D0BWP7T port map(A1 => n_203, A2 => n_995, B => n_1005, C => n_455, ZN => n_1026);
  g29187 : OAI211D0BWP7T port map(A1 => n_203, A2 => n_987, B => n_1004, C => n_459, ZN => n_1025);
  g29188 : INR4D0BWP7T port map(A1 => n_999, B1 => corner_count(8), B2 => corner_count(9), B3 => corner_count(10), ZN => n_1024);
  g29189 : OAI211D0BWP7T port map(A1 => n_203, A2 => n_984, B => n_1006, C => n_447, ZN => n_1023);
  g29190 : MOAI22D0BWP7T port map(A1 => n_1008, A2 => new_tail(5), B1 => n_1008, B2 => new_tail(5), ZN => n_1022);
  g29191 : MOAI22D0BWP7T port map(A1 => n_1014, A2 => new_tail(3), B1 => n_1014, B2 => new_tail(3), ZN => n_1021);
  g29192 : MOAI22D0BWP7T port map(A1 => n_1011, A2 => new_tail(1), B1 => n_1011, B2 => new_tail(1), ZN => n_1020);
  g29193 : ND2D0BWP7T port map(A1 => n_1015, A2 => new_tail(4), ZN => n_1019);
  g29194 : OAI211D0BWP7T port map(A1 => n_205, A2 => n_994, B => n_998, C => n_443, ZN => n_1018);
  g29195 : OAI221D0BWP7T port map(A1 => n_985, A2 => n_203, B1 => n_155, B2 => n_208, C => n_1009, ZN => n_1017);
  g29196 : OAI221D0BWP7T port map(A1 => n_997, A2 => n_203, B1 => n_155, B2 => n_206, C => n_1010, ZN => n_1016);
  g29197 : OA21D0BWP7T port map(A1 => n_985, A2 => n_205, B => n_453, Z => n_1010);
  g29198 : OA21D0BWP7T port map(A1 => n_997, A2 => n_205, B => n_445, Z => n_1009);
  g29199 : AN4D1BWP7T port map(A1 => n_977, A2 => n_786, A3 => n_787, A4 => n_743, Z => n_1015);
  g29200 : AN4D1BWP7T port map(A1 => n_978, A2 => n_783, A3 => n_784, A4 => n_744, Z => n_1014);
  g29201 : AN4D1BWP7T port map(A1 => n_979, A2 => n_780, A3 => n_781, A4 => n_745, Z => n_1013);
  g29202 : AN4D1BWP7T port map(A1 => n_980, A2 => n_777, A3 => n_778, A4 => n_746, Z => n_1012);
  g29203 : AN4D1BWP7T port map(A1 => n_981, A2 => n_774, A3 => n_775, A4 => n_747, Z => n_1011);
  g29204 : AOI22D0BWP7T port map(A1 => n_996, A2 => n_202, B1 => n_1737, B2 => head(1), ZN => n_1007);
  g29205 : AOI22D0BWP7T port map(A1 => n_983, A2 => n_204, B1 => n_1737, B2 => head(3), ZN => n_1006);
  g29206 : AOI22D0BWP7T port map(A1 => n_996, A2 => n_204, B1 => n_1737, B2 => head(6), ZN => n_1005);
  g29207 : AOI22D0BWP7T port map(A1 => n_986, A2 => n_204, B1 => n_1737, B2 => head(9), ZN => n_1004);
  g29208 : AOI22D0BWP7T port map(A1 => n_983, A2 => n_202, B1 => n_1737, B2 => head(8), ZN => n_1003);
  g29209 : AOI22D0BWP7T port map(A1 => n_986, A2 => n_202, B1 => n_1737, B2 => head(4), ZN => n_1002);
  g29210 : MAOI22D0BWP7T port map(A1 => n_1737, A2 => head(5), B1 => n_994, B2 => n_203, ZN => n_1001);
  g29211 : AN4D1BWP7T port map(A1 => n_982, A2 => n_790, A3 => n_791, A4 => n_717, Z => n_1008);
  g29216 : AOI21D0BWP7T port map(A1 => n_1735, A2 => snake_output1(5), B => n_993, ZN => n_1000);
  g29217 : INR4D0BWP7T port map(A1 => n_969, B1 => corner_count(5), B2 => corner_count(6), B3 => corner_count(7), ZN => n_999);
  g29219 : MAOI22D0BWP7T port map(A1 => n_1737, A2 => head(0), B1 => n_976, B2 => n_203, ZN => n_998);
  g29220 : OAI21D0BWP7T port map(A1 => n_599, A2 => n_230, B => n_975, ZN => n_993);
  g29221 : ND4D0BWP7T port map(A1 => n_966, A2 => n_818, A3 => n_819, A4 => n_730, ZN => n_992);
  g29222 : ND4D0BWP7T port map(A1 => n_965, A2 => n_815, A3 => n_816, A4 => n_729, ZN => n_991);
  g29223 : ND4D0BWP7T port map(A1 => n_964, A2 => n_813, A3 => n_820, A4 => n_726, ZN => n_990);
  g29224 : ND4D0BWP7T port map(A1 => n_957, A2 => n_828, A3 => n_827, A4 => n_724, ZN => n_989);
  g29225 : ND4D0BWP7T port map(A1 => n_962, A2 => n_831, A3 => n_830, A4 => n_722, ZN => n_988);
  g29226 : AN4D1BWP7T port map(A1 => n_958, A2 => n_711, A3 => n_654, A4 => n_655, Z => n_997);
  g29227 : ND4D0BWP7T port map(A1 => n_959, A2 => n_713, A3 => n_586, A4 => n_658, ZN => n_996);
  g29228 : AN4D1BWP7T port map(A1 => n_960, A2 => n_715, A3 => n_665, A4 => n_666, Z => n_995);
  g29229 : AN4D1BWP7T port map(A1 => n_961, A2 => n_720, A3 => n_624, A4 => n_678, Z => n_994);
  g29230 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(5), B1 => n_605, B2 => snake_output21(5), C => n_972, ZN => n_982);
  g29231 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(1), B1 => n_605, B2 => snake_output21(1), C => n_967, ZN => n_981);
  g29232 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(2), B1 => n_605, B2 => snake_output21(2), C => n_968, ZN => n_980);
  g29233 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(0), B1 => n_605, B2 => snake_output21(0), C => n_974, ZN => n_979);
  g29234 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(3), B1 => n_605, B2 => snake_output21(3), C => n_970, ZN => n_978);
  g29235 : AOI221D0BWP7T port map(A1 => n_0, A2 => snake_output16(4), B1 => n_605, B2 => snake_output21(4), C => n_971, ZN => n_977);
  g29236 : AN4D1BWP7T port map(A1 => n_954, A2 => n_705, A3 => n_638, A4 => n_639, Z => n_987);
  g29237 : ND4D0BWP7T port map(A1 => n_953, A2 => n_704, A3 => n_576, A4 => n_634, ZN => n_986);
  g29238 : AN4D1BWP7T port map(A1 => n_963, A2 => n_710, A3 => n_582, A4 => n_649, Z => n_985);
  g29239 : AN4D1BWP7T port map(A1 => n_955, A2 => n_707, A3 => n_579, A4 => n_642, Z => n_984);
  g29240 : ND4D0BWP7T port map(A1 => n_956, A2 => n_708, A3 => n_645, A4 => n_646, ZN => n_983);
  g29242 : AOI31D0BWP7T port map(A1 => n_427, A2 => n_226, A3 => snake_output13(5), B => n_973, ZN => n_975);
  g29243 : AN4D1BWP7T port map(A1 => n_951, A2 => n_719, A3 => n_589, A4 => n_668, Z => n_976);
  g29244 : ND4D0BWP7T port map(A1 => n_947, A2 => n_735, A3 => n_568, A4 => n_567, ZN => n_974);
  g29245 : IOA21D0BWP7T port map(A1 => n_940, A2 => n_1736, B => n_822, ZN => n_973);
  g29246 : ND4D0BWP7T port map(A1 => n_950, A2 => n_731, A3 => n_574, A4 => n_573, ZN => n_972);
  g29247 : ND4D0BWP7T port map(A1 => n_949, A2 => n_732, A3 => n_571, A4 => n_572, ZN => n_971);
  g29248 : ND4D0BWP7T port map(A1 => n_948, A2 => n_733, A3 => n_569, A4 => n_570, ZN => n_970);
  g29249 : INR4D0BWP7T port map(A1 => n_927, B1 => corner_count(19), B2 => corner_count(17), B3 => corner_count(18), ZN => n_969);
  g29250 : ND4D0BWP7T port map(A1 => n_946, A2 => n_736, A3 => n_591, A4 => n_578, ZN => n_968);
  g29251 : ND4D0BWP7T port map(A1 => n_945, A2 => n_737, A3 => n_593, A4 => n_592, ZN => n_967);
  g29252 : AOI221D0BWP7T port map(A1 => n_465, A2 => snake_output15(0), B1 => n_560, B2 => snake_output21(0), C => n_944, ZN => n_966);
  g29253 : AOI221D0BWP7T port map(A1 => n_465, A2 => snake_output15(1), B1 => n_560, B2 => snake_output21(1), C => n_943, ZN => n_965);
  g29254 : AOI221D0BWP7T port map(A1 => n_465, A2 => snake_output15(2), B1 => n_560, B2 => snake_output21(2), C => n_942, ZN => n_964);
  g29255 : AOI221D0BWP7T port map(A1 => n_562, A2 => snake_output23(2), B1 => n_534, B2 => snake_output18(2), C => n_938, ZN => n_963);
  g29256 : AOI221D0BWP7T port map(A1 => n_465, A2 => snake_output15(4), B1 => n_560, B2 => snake_output21(4), C => n_935, ZN => n_962);
  g29257 : AOI221D0BWP7T port map(A1 => n_515, A2 => snake_output17(0), B1 => n_602, B2 => snake_output22(0), C => n_934, ZN => n_961);
  g29258 : AOI221D0BWP7T port map(A1 => n_515, A2 => snake_output17(1), B1 => n_602, B2 => snake_output22(1), C => n_933, ZN => n_960);
  g29259 : AOI221D0BWP7T port map(A1 => n_562, A2 => snake_output23(1), B1 => n_534, B2 => snake_output18(1), C => n_939, ZN => n_959);
  g29260 : AOI221D0BWP7T port map(A1 => n_515, A2 => snake_output17(2), B1 => n_602, B2 => snake_output22(2), C => n_932, ZN => n_958);
  g29261 : AOI221D0BWP7T port map(A1 => n_465, A2 => snake_output15(3), B1 => n_560, B2 => snake_output21(3), C => n_941, ZN => n_957);
  g29262 : AOI221D0BWP7T port map(A1 => n_515, A2 => snake_output17(3), B1 => n_602, B2 => snake_output22(3), C => n_931, ZN => n_956);
  g29263 : AOI221D0BWP7T port map(A1 => n_562, A2 => snake_output23(3), B1 => n_534, B2 => snake_output18(3), C => n_937, ZN => n_955);
  g29264 : AOI221D0BWP7T port map(A1 => n_515, A2 => snake_output17(4), B1 => n_602, B2 => snake_output22(4), C => n_930, ZN => n_954);
  g29265 : AOI221D0BWP7T port map(A1 => n_562, A2 => snake_output23(4), B1 => n_534, B2 => snake_output18(4), C => n_936, ZN => n_953);
  g29266 : AO22D0BWP7T port map(A1 => n_940, A2 => n_192, B1 => snake_output0(5), B2 => n_1737, Z => n_952);
  g29267 : AOI221D0BWP7T port map(A1 => n_562, A2 => snake_output23(0), B1 => n_534, B2 => snake_output18(0), C => n_922, ZN => n_951);
  g29268 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(5), B1 => n_518, B2 => snake_output15(5), C => n_928, ZN => n_950);
  g29269 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(4), B1 => n_518, B2 => snake_output15(4), C => n_929, ZN => n_949);
  g29270 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(3), B1 => n_518, B2 => snake_output15(3), C => n_926, ZN => n_948);
  g29271 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(0), B1 => n_518, B2 => snake_output15(0), C => n_923, ZN => n_947);
  g29272 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(2), B1 => n_518, B2 => snake_output15(2), C => n_924, ZN => n_946);
  g29273 : AOI221D0BWP7T port map(A1 => n_517, A2 => snake_output14(1), B1 => n_518, B2 => snake_output15(1), C => n_925, ZN => n_945);
  g29274 : ND4D0BWP7T port map(A1 => n_906, A2 => n_861, A3 => n_853, A4 => n_680, ZN => n_944);
  g29275 : ND4D0BWP7T port map(A1 => n_910, A2 => n_826, A3 => n_728, A4 => n_814, ZN => n_943);
  g29276 : ND4D0BWP7T port map(A1 => n_909, A2 => n_825, A3 => n_852, A4 => n_821, ZN => n_942);
  g29277 : ND4D0BWP7T port map(A1 => n_908, A2 => n_824, A3 => n_851, A4 => n_829, ZN => n_941);
  g29278 : ND4D0BWP7T port map(A1 => n_916, A2 => n_712, A3 => n_657, A4 => n_628, ZN => n_939);
  g29279 : ND4D0BWP7T port map(A1 => n_915, A2 => n_709, A3 => n_648, A4 => n_627, ZN => n_938);
  g29280 : ND4D0BWP7T port map(A1 => n_914, A2 => n_706, A3 => n_641, A4 => n_626, ZN => n_937);
  g29281 : ND4D0BWP7T port map(A1 => n_913, A2 => n_703, A3 => n_633, A4 => n_625, ZN => n_936);
  g29282 : ND4D0BWP7T port map(A1 => n_907, A2 => n_823, A3 => n_850, A4 => n_832, ZN => n_935);
  g29283 : ND4D0BWP7T port map(A1 => n_921, A2 => n_671, A3 => n_833, A4 => n_834, ZN => n_934);
  g29284 : ND4D0BWP7T port map(A1 => n_920, A2 => n_663, A3 => n_838, A4 => n_839, ZN => n_933);
  g29285 : ND4D0BWP7T port map(A1 => n_919, A2 => n_653, A3 => n_806, A4 => n_805, ZN => n_932);
  g29286 : ND4D0BWP7T port map(A1 => n_918, A2 => n_644, A3 => n_801, A4 => n_800, ZN => n_931);
  g29287 : ND4D0BWP7T port map(A1 => n_917, A2 => n_637, A3 => n_796, A4 => n_795, ZN => n_930);
  g29288 : ND4D0BWP7T port map(A1 => n_912, A2 => n_718, A3 => n_716, A4 => n_672, ZN => n_940);
  g29289 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(4), B => n_911, Z => n_929);
  g29290 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(5), B => n_901, Z => n_928);
  g29291 : INR4D0BWP7T port map(A1 => n_885, B1 => corner_count(22), B2 => corner_count(21), B3 => corner_count(20), ZN => n_927);
  g29292 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(3), B => n_905, Z => n_926);
  g29293 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(1), B => n_902, Z => n_925);
  g29294 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(2), B => n_903, Z => n_924);
  g29295 : AO21D0BWP7T port map(A1 => n_604, A2 => snake_output24(0), B => n_904, Z => n_923);
  g29296 : ND4D0BWP7T port map(A1 => n_898, A2 => n_837, A3 => n_836, A4 => n_588, ZN => n_922);
  g29297 : AOI221D0BWP7T port map(A1 => n_498, A2 => snake_output3(0), B1 => n_510, B2 => snake_output2(0), C => n_899, ZN => n_921);
  g29298 : AOI221D0BWP7T port map(A1 => n_498, A2 => snake_output3(1), B1 => n_510, B2 => snake_output2(1), C => n_900, ZN => n_920);
  g29299 : AOI221D0BWP7T port map(A1 => n_498, A2 => snake_output3(2), B1 => n_510, B2 => snake_output2(2), C => n_896, ZN => n_919);
  g29300 : AOI221D0BWP7T port map(A1 => n_498, A2 => snake_output3(3), B1 => n_510, B2 => snake_output2(3), C => n_894, ZN => n_918);
  g29301 : AOI221D0BWP7T port map(A1 => n_498, A2 => snake_output3(4), B1 => n_510, B2 => snake_output2(4), C => n_892, ZN => n_917);
  g29302 : AOI221D0BWP7T port map(A1 => n_475, A2 => snake_output14(1), B1 => n_418, B2 => snake_output13(1), C => n_897, ZN => n_916);
  g29303 : AOI221D0BWP7T port map(A1 => n_514, A2 => snake_output11(2), B1 => n_475, B2 => snake_output14(2), C => n_893, ZN => n_915);
  g29304 : AOI221D0BWP7T port map(A1 => n_514, A2 => snake_output11(3), B1 => n_475, B2 => snake_output14(3), C => n_895, ZN => n_914);
  g29305 : AOI221D0BWP7T port map(A1 => n_514, A2 => snake_output11(4), B1 => n_475, B2 => snake_output14(4), C => n_891, ZN => n_913);
  g29306 : NR3D0BWP7T port map(A1 => n_869, A2 => n_871, A3 => n_810, ZN => n_912);
  g29307 : ND4D0BWP7T port map(A1 => n_877, A2 => n_848, A3 => n_785, A4 => n_772, ZN => n_911);
  g29308 : AOI221D0BWP7T port map(A1 => n_752, A2 => snake_output8(1), B1 => n_480, B2 => snake_output22(1), C => n_883, ZN => n_910);
  g29309 : AOI221D0BWP7T port map(A1 => n_618, A2 => snake_output10(2), B1 => n_480, B2 => snake_output22(2), C => n_882, ZN => n_909);
  g29310 : AOI221D0BWP7T port map(A1 => n_618, A2 => snake_output10(3), B1 => n_480, B2 => snake_output22(3), C => n_881, ZN => n_908);
  g29311 : AOI221D0BWP7T port map(A1 => n_618, A2 => snake_output10(4), B1 => n_480, B2 => snake_output22(4), C => n_880, ZN => n_907);
  g29312 : AOI221D0BWP7T port map(A1 => n_618, A2 => snake_output10(0), B1 => n_480, B2 => snake_output22(0), C => n_884, ZN => n_906);
  g29313 : ND4D0BWP7T port map(A1 => n_876, A2 => n_847, A3 => n_782, A4 => n_771, ZN => n_905);
  g29314 : ND4D0BWP7T port map(A1 => n_875, A2 => n_846, A3 => n_779, A4 => n_770, ZN => n_904);
  g29315 : ND4D0BWP7T port map(A1 => n_874, A2 => n_845, A3 => n_776, A4 => n_769, ZN => n_903);
  g29316 : ND4D0BWP7T port map(A1 => n_873, A2 => n_844, A3 => n_773, A4 => n_768, ZN => n_902);
  g29317 : ND4D0BWP7T port map(A1 => n_878, A2 => n_849, A3 => n_788, A4 => n_789, ZN => n_901);
  g29318 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(1), B => n_870, Z => n_900);
  g29319 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(0), B => n_872, Z => n_899);
  g29320 : AOI221D0BWP7T port map(A1 => n_510, A2 => snake_output1(0), B1 => n_532, B2 => snake_output5(0), C => n_879, ZN => n_898);
  g29321 : AO21D0BWP7T port map(A1 => n_621, A2 => snake_output24(1), B => n_868, Z => n_897);
  g29322 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(2), B => n_867, Z => n_896);
  g29323 : AO21D0BWP7T port map(A1 => n_621, A2 => snake_output24(3), B => n_864, Z => n_895);
  g29324 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(3), B => n_865, Z => n_894);
  g29325 : AO21D0BWP7T port map(A1 => n_621, A2 => snake_output24(2), B => n_866, Z => n_893);
  g29326 : AO21D0BWP7T port map(A1 => n_611, A2 => snake_output24(4), B => n_863, Z => n_892);
  g29327 : AO21D0BWP7T port map(A1 => n_621, A2 => snake_output24(4), B => n_862, Z => n_891);
  g29355 : INR4D0BWP7T port map(A1 => n_734, B1 => corner_count(25), B2 => corner_count(24), B3 => corner_count(23), ZN => n_885);
  g29356 : ND3D0BWP7T port map(A1 => n_843, A2 => n_738, A3 => n_681, ZN => n_884);
  g29357 : ND3D0BWP7T port map(A1 => n_857, A2 => n_739, A3 => n_682, ZN => n_883);
  g29358 : ND3D0BWP7T port map(A1 => n_856, A2 => n_740, A3 => n_683, ZN => n_882);
  g29359 : ND3D0BWP7T port map(A1 => n_855, A2 => n_741, A3 => n_677, ZN => n_881);
  g29360 : ND3D0BWP7T port map(A1 => n_854, A2 => n_742, A3 => n_675, ZN => n_880);
  g29361 : AO21D0BWP7T port map(A1 => n_621, A2 => snake_output24(0), B => n_858, Z => n_879);
  g29362 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(5), B1 => n_841, B2 => snake_output7(5), ZN => n_878);
  g29363 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(4), B1 => n_841, B2 => snake_output7(4), ZN => n_877);
  g29364 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(3), B1 => n_841, B2 => snake_output7(3), ZN => n_876);
  g29365 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(0), B1 => n_841, B2 => snake_output7(0), ZN => n_875);
  g29366 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(2), B1 => n_841, B2 => snake_output7(2), ZN => n_874);
  g29367 : AOI22D0BWP7T port map(A1 => n_842, A2 => snake_output6(1), B1 => n_841, B2 => snake_output7(1), ZN => n_873);
  g29368 : ND4D0BWP7T port map(A1 => n_835, A2 => n_670, A3 => n_669, A4 => n_590, ZN => n_872);
  g29369 : ND4D0BWP7T port map(A1 => n_808, A2 => n_662, A3 => n_660, A4 => n_714, ZN => n_871);
  g29370 : ND4D0BWP7T port map(A1 => n_840, A2 => n_661, A3 => n_659, A4 => n_587, ZN => n_870);
  g29371 : ND4D0BWP7T port map(A1 => n_652, A2 => n_584, A3 => n_807, A4 => n_630, ZN => n_869);
  g29372 : ND4D0BWP7T port map(A1 => n_809, A2 => n_767, A3 => n_585, A4 => n_656, ZN => n_868);
  g29373 : ND4D0BWP7T port map(A1 => n_804, A2 => n_651, A3 => n_650, A4 => n_583, ZN => n_867);
  g29374 : ND4D0BWP7T port map(A1 => n_803, A2 => n_802, A3 => n_581, A4 => n_647, ZN => n_866);
  g29375 : ND4D0BWP7T port map(A1 => n_799, A2 => n_632, A3 => n_643, A4 => n_580, ZN => n_865);
  g29376 : ND4D0BWP7T port map(A1 => n_797, A2 => n_594, A3 => n_798, A4 => n_640, ZN => n_864);
  g29377 : ND4D0BWP7T port map(A1 => n_794, A2 => n_636, A3 => n_635, A4 => n_577, ZN => n_863);
  g29378 : ND4D0BWP7T port map(A1 => n_792, A2 => n_793, A3 => n_575, A4 => n_631, ZN => n_862);
  g29382 : AOI221D0BWP7T port map(A1 => n_538, A2 => snake_output16(0), B1 => n_558, B2 => snake_output13(0), C => n_817, ZN => n_861);
  g29395 : OAI21D0BWP7T port map(A1 => n_1, A2 => n_1701, B => n_195, ZN => n_890);
  g29396 : AOI21D0BWP7T port map(A1 => n_754, A2 => n_222, B => n_194, ZN => n_886);
  g29397 : AOI21D0BWP7T port map(A1 => n_754, A2 => n_212, B => n_194, ZN => n_887);
  g29398 : OAI21D0BWP7T port map(A1 => n_753, A2 => n_217, B => n_195, ZN => n_889);
  g29399 : ND4D0BWP7T port map(A1 => n_748, A2 => n_667, A3 => n_629, A4 => n_527, ZN => n_858);
  g29400 : AOI222D0BWP7T port map(A1 => n_614, A2 => snake_output1(1), B1 => n_616, B2 => snake_output14(1), C1 => n_751, C2 => snake_output5(1), ZN => n_857);
  g29401 : AOI222D0BWP7T port map(A1 => n_614, A2 => snake_output1(2), B1 => n_616, B2 => snake_output14(2), C1 => n_751, C2 => snake_output5(2), ZN => n_856);
  g29402 : AOI222D0BWP7T port map(A1 => n_614, A2 => snake_output1(3), B1 => n_616, B2 => snake_output14(3), C1 => n_751, C2 => snake_output5(3), ZN => n_855);
  g29403 : AOI222D0BWP7T port map(A1 => n_614, A2 => snake_output1(4), B1 => n_616, B2 => snake_output14(4), C1 => n_751, C2 => snake_output5(4), ZN => n_854);
  g29404 : AOI22D0BWP7T port map(A1 => n_752, A2 => snake_output8(0), B1 => n_615, B2 => snake_output7(0), ZN => n_853);
  g29405 : AOI22D0BWP7T port map(A1 => n_752, A2 => snake_output8(2), B1 => n_557, B2 => snake_output11(2), ZN => n_852);
  g29406 : AOI22D0BWP7T port map(A1 => n_752, A2 => snake_output8(3), B1 => n_557, B2 => snake_output11(3), ZN => n_851);
  g29407 : AOI22D0BWP7T port map(A1 => n_752, A2 => snake_output8(4), B1 => n_557, B2 => snake_output11(4), ZN => n_850);
  g29408 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(5), B1 => n_749, B2 => snake_output3(5), ZN => n_849);
  g29409 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(4), B1 => n_749, B2 => snake_output3(4), ZN => n_848);
  g29410 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(3), B1 => n_749, B2 => snake_output3(3), ZN => n_847);
  g29411 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(0), B1 => n_749, B2 => snake_output3(0), ZN => n_846);
  g29412 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(2), B1 => n_749, B2 => snake_output3(2), ZN => n_845);
  g29413 : AOI22D0BWP7T port map(A1 => n_750, A2 => snake_output2(1), B1 => n_749, B2 => snake_output3(1), ZN => n_844);
  g29414 : AOI222D0BWP7T port map(A1 => n_614, A2 => snake_output1(0), B1 => n_616, B2 => snake_output14(0), C1 => n_751, C2 => snake_output5(0), ZN => n_843);
  g29415 : OAI21D0BWP7T port map(A1 => n_753, A2 => n_220, B => n_195, ZN => n_888);
  g29416 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output8(1), B1 => n_554, B2 => snake_output9(1), ZN => n_840);
  g29417 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output4(1), B1 => n_500, B2 => snake_output5(1), ZN => n_839);
  g29418 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(1), B1 => n_532, B2 => snake_output6(1), ZN => n_838);
  g29419 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output7(0), B1 => n_685, B2 => snake_output6(0), ZN => n_837);
  g29420 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output3(0), B1 => n_498, B2 => snake_output2(0), ZN => n_836);
  g29421 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output8(0), B1 => n_554, B2 => snake_output9(0), ZN => n_835);
  g29422 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output4(0), B1 => n_500, B2 => snake_output5(0), ZN => n_834);
  g29423 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(0), B1 => n_532, B2 => snake_output6(0), ZN => n_833);
  g29424 : AOI22D0BWP7T port map(A1 => n_698, A2 => snake_output9(4), B1 => n_613, B2 => snake_output12(4), ZN => n_832);
  g29425 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(4), B1 => n_697, B2 => snake_output23(4), ZN => n_831);
  g29426 : AOI22D0BWP7T port map(A1 => n_695, A2 => snake_output19(4), B1 => n_696, B2 => snake_output24(4), ZN => n_830);
  g29427 : AOI22D0BWP7T port map(A1 => n_698, A2 => snake_output9(3), B1 => n_613, B2 => snake_output12(3), ZN => n_829);
  g29428 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(3), B1 => n_697, B2 => snake_output23(3), ZN => n_828);
  g29429 : AOI22D0BWP7T port map(A1 => n_695, A2 => snake_output19(3), B1 => n_696, B2 => snake_output24(3), ZN => n_827);
  g29430 : AOI221D0BWP7T port map(A1 => n_561, A2 => snake_output6(1), B1 => n_558, B2 => snake_output13(1), C => n_727, ZN => n_826);
  g29431 : AOI221D0BWP7T port map(A1 => n_561, A2 => snake_output6(2), B1 => n_558, B2 => snake_output13(2), C => n_725, ZN => n_825);
  g29432 : AOI221D0BWP7T port map(A1 => n_561, A2 => snake_output6(3), B1 => n_558, B2 => snake_output13(3), C => n_723, ZN => n_824);
  g29433 : AOI221D0BWP7T port map(A1 => n_561, A2 => snake_output6(4), B1 => n_558, B2 => snake_output13(4), C => n_721, ZN => n_823);
  g29434 : OAI31D0BWP7T port map(A1 => n_600, A2 => n_1732, A3 => n_1737, B => snake_output0(5), ZN => n_822);
  g29435 : AOI22D0BWP7T port map(A1 => n_698, A2 => snake_output9(2), B1 => n_613, B2 => snake_output12(2), ZN => n_821);
  g29436 : AOI22D0BWP7T port map(A1 => n_695, A2 => snake_output19(2), B1 => n_696, B2 => snake_output24(2), ZN => n_820);
  g29437 : AOI22D0BWP7T port map(A1 => n_695, A2 => snake_output19(0), B1 => n_696, B2 => snake_output24(0), ZN => n_819);
  g29438 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(0), B1 => n_697, B2 => snake_output23(0), ZN => n_818);
  g29439 : AO22D0BWP7T port map(A1 => n_698, A2 => snake_output9(0), B1 => snake_output12(0), B2 => n_613, Z => n_817);
  g29440 : AOI22D0BWP7T port map(A1 => n_695, A2 => snake_output19(1), B1 => n_696, B2 => snake_output24(1), ZN => n_816);
  g29441 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(1), B1 => n_697, B2 => snake_output23(1), ZN => n_815);
  g29442 : AOI22D0BWP7T port map(A1 => n_698, A2 => snake_output9(1), B1 => n_618, B2 => snake_output10(1), ZN => n_814);
  g29443 : AOI22D0BWP7T port map(A1 => n_620, A2 => snake_output17(2), B1 => n_697, B2 => snake_output23(2), ZN => n_813);
  g29446 : NR2D0BWP7T port map(A1 => n_755, A2 => corner_count(0), ZN => n_842);
  g29447 : NR2D0BWP7T port map(A1 => n_755, A2 => n_146, ZN => n_841);
  g29457 : AOI21D1BWP7T port map(A1 => n_700, A2 => n_1700, B => n_194, ZN => n_860);
  g29459 : OAI21D0BWP7T port map(A1 => n_701, A2 => n_1700, B => n_195, ZN => n_859);
  g29460 : MOAI22D0BWP7T port map(A1 => n_664, A2 => n_477, B1 => n_515, B2 => snake_output18(5), ZN => n_810);
  g29461 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output7(1), B1 => n_685, B2 => snake_output6(1), ZN => n_809);
  g29462 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output8(5), B1 => n_554, B2 => snake_output10(5), ZN => n_808);
  g29463 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output5(5), B1 => n_496, B2 => snake_output2(5), ZN => n_807);
  g29464 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(2), B1 => n_532, B2 => snake_output6(2), ZN => n_806);
  g29465 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output4(2), B1 => n_500, B2 => snake_output5(2), ZN => n_805);
  g29466 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output8(2), B1 => n_554, B2 => snake_output9(2), ZN => n_804);
  g29467 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output7(2), B1 => n_685, B2 => snake_output6(2), ZN => n_803);
  g29468 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output3(2), B1 => n_498, B2 => snake_output2(2), ZN => n_802);
  g29469 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(3), B1 => n_532, B2 => snake_output6(3), ZN => n_801);
  g29470 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output4(3), B1 => n_500, B2 => snake_output5(3), ZN => n_800);
  g29471 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output8(3), B1 => n_554, B2 => snake_output9(3), ZN => n_799);
  g29472 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output3(3), B1 => n_496, B2 => snake_output0(3), ZN => n_798);
  g29473 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output7(3), B1 => n_685, B2 => snake_output6(3), ZN => n_797);
  g29474 : AOI22D0BWP7T port map(A1 => n_685, A2 => snake_output7(4), B1 => n_532, B2 => snake_output6(4), ZN => n_796);
  g29475 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output4(4), B1 => n_500, B2 => snake_output5(4), ZN => n_795);
  g29476 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output8(4), B1 => n_554, B2 => snake_output9(4), ZN => n_794);
  g29477 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output3(4), B1 => n_498, B2 => snake_output2(4), ZN => n_793);
  g29478 : AOI22D0BWP7T port map(A1 => n_688, A2 => snake_output7(4), B1 => n_685, B2 => snake_output6(4), ZN => n_792);
  g29479 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(5), B1 => n_606, B2 => snake_output18(5), ZN => n_791);
  g29480 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(5), B1 => n_608, B2 => snake_output17(5), ZN => n_790);
  g29481 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(5), B1 => n_693, B2 => snake_output5(5), ZN => n_789);
  g29482 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(5), B1 => n_689, B2 => snake_output1(5), ZN => n_788);
  g29483 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(4), B1 => n_606, B2 => snake_output18(4), ZN => n_787);
  g29484 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(4), B1 => n_608, B2 => snake_output17(4), ZN => n_786);
  g29485 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(4), B1 => n_689, B2 => snake_output1(4), ZN => n_785);
  g29486 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(3), B1 => n_606, B2 => snake_output18(3), ZN => n_784);
  g29487 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(3), B1 => n_608, B2 => snake_output17(3), ZN => n_783);
  g29488 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(3), B1 => n_689, B2 => snake_output1(3), ZN => n_782);
  g29489 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(0), B1 => n_606, B2 => snake_output18(0), ZN => n_781);
  g29490 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(0), B1 => n_608, B2 => snake_output17(0), ZN => n_780);
  g29491 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(0), B1 => n_689, B2 => snake_output1(0), ZN => n_779);
  g29492 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(2), B1 => n_606, B2 => snake_output18(2), ZN => n_778);
  g29493 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(2), B1 => n_608, B2 => snake_output17(2), ZN => n_777);
  g29494 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(2), B1 => n_689, B2 => snake_output1(2), ZN => n_776);
  g29495 : AOI22D0BWP7T port map(A1 => n_692, A2 => snake_output22(1), B1 => n_606, B2 => snake_output18(1), ZN => n_775);
  g29496 : AOI22D0BWP7T port map(A1 => n_691, A2 => snake_output23(1), B1 => n_608, B2 => snake_output17(1), ZN => n_774);
  g29497 : AOI22D0BWP7T port map(A1 => n_694, A2 => snake_output0(1), B1 => n_689, B2 => snake_output1(1), ZN => n_773);
  g29498 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(4), B1 => n_693, B2 => snake_output5(4), ZN => n_772);
  g29499 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(3), B1 => n_693, B2 => snake_output5(3), ZN => n_771);
  g29500 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(0), B1 => n_693, B2 => snake_output5(0), ZN => n_770);
  g29501 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(2), B1 => n_693, B2 => snake_output5(2), ZN => n_769);
  g29502 : AOI22D0BWP7T port map(A1 => n_690, A2 => snake_output4(1), B1 => n_693, B2 => snake_output5(1), ZN => n_768);
  g29503 : AOI22D0BWP7T port map(A1 => n_687, A2 => snake_output3(1), B1 => n_498, B2 => snake_output2(1), ZN => n_767);
  g29567 : CKND1BWP7T port map(I => n_754, ZN => n_753);
  g29568 : AOI22D0BWP7T port map(A1 => n_617, A2 => snake_output8(0), B1 => n_512, B2 => snake_output9(0), ZN => n_748);
  g29569 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(1), B1 => n_609, B2 => snake_output20(1), ZN => n_747);
  g29570 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(2), B1 => n_609, B2 => snake_output20(2), ZN => n_746);
  g29571 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(0), B1 => n_609, B2 => snake_output20(0), ZN => n_745);
  g29572 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(3), B1 => n_609, B2 => snake_output20(3), ZN => n_744);
  g29573 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(4), B1 => n_609, B2 => snake_output20(4), ZN => n_743);
  g29574 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(4), B1 => n_537, B2 => snake_output2(4), ZN => n_742);
  g29575 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(3), B1 => n_537, B2 => snake_output2(3), ZN => n_741);
  g29576 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(2), B1 => n_537, B2 => snake_output2(2), ZN => n_740);
  g29577 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(1), B1 => n_537, B2 => snake_output2(1), ZN => n_739);
  g29578 : AOI22D0BWP7T port map(A1 => n_597, A2 => snake_output0(0), B1 => n_537, B2 => snake_output2(0), ZN => n_738);
  g29579 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(1), B1 => n_516, B2 => snake_output9(1), ZN => n_737);
  g29580 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(2), B1 => n_516, B2 => snake_output9(2), ZN => n_736);
  g29581 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(0), B1 => n_516, B2 => snake_output9(0), ZN => n_735);
  g29582 : INR4D0BWP7T port map(A1 => n_528, B1 => corner_count(28), B2 => corner_count(27), B3 => corner_count(26), ZN => n_734);
  g29583 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(3), B1 => n_516, B2 => snake_output9(3), ZN => n_733);
  g29585 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(4), B1 => n_516, B2 => snake_output9(4), ZN => n_732);
  g29586 : AOI22D0BWP7T port map(A1 => n_603, A2 => snake_output8(5), B1 => n_516, B2 => snake_output9(5), ZN => n_731);
  g29587 : AOI22D0BWP7T port map(A1 => n_612, A2 => snake_output20(0), B1 => n_556, B2 => snake_output18(0), ZN => n_730);
  g29588 : AOI22D0BWP7T port map(A1 => n_612, A2 => snake_output20(1), B1 => n_556, B2 => snake_output18(1), ZN => n_729);
  g29589 : AOI22D0BWP7T port map(A1 => n_557, A2 => snake_output11(1), B1 => n_613, B2 => snake_output12(1), ZN => n_728);
  g29590 : AO22D0BWP7T port map(A1 => n_538, A2 => snake_output16(1), B1 => snake_output7(1), B2 => n_615, Z => n_727);
  g29591 : AOI22D0BWP7T port map(A1 => n_612, A2 => snake_output20(2), B1 => n_556, B2 => snake_output18(2), ZN => n_726);
  g29592 : AO22D0BWP7T port map(A1 => n_538, A2 => snake_output16(2), B1 => snake_output7(2), B2 => n_615, Z => n_725);
  g29593 : AOI22D0BWP7T port map(A1 => n_612, A2 => snake_output20(3), B1 => n_556, B2 => snake_output18(3), ZN => n_724);
  g29594 : AO22D0BWP7T port map(A1 => n_538, A2 => snake_output16(3), B1 => snake_output7(3), B2 => n_615, Z => n_723);
  g29595 : AOI22D0BWP7T port map(A1 => n_612, A2 => snake_output20(4), B1 => n_556, B2 => snake_output18(4), ZN => n_722);
  g29596 : AO22D0BWP7T port map(A1 => n_538, A2 => snake_output16(4), B1 => snake_output7(4), B2 => n_615, Z => n_721);
  g29597 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output18(0), B1 => n_502, B2 => snake_output20(0), ZN => n_720);
  g29598 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output17(0), B1 => n_602, B2 => snake_output21(0), ZN => n_719);
  g29599 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output19(5), B1 => n_534, B2 => snake_output20(5), ZN => n_718);
  g29600 : AOI22D0BWP7T port map(A1 => n_607, A2 => snake_output19(5), B1 => n_609, B2 => snake_output20(5), ZN => n_717);
  g29601 : AOI22D0BWP7T port map(A1 => n_602, A2 => n_1053, B1 => n_502, B2 => snake_output21(5), ZN => n_716);
  g29602 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output18(1), B1 => n_502, B2 => snake_output20(1), ZN => n_715);
  g29603 : AOI22D0BWP7T port map(A1 => n_622, A2 => snake_output9(5), B1 => n_512, B2 => snake_output11(5), ZN => n_714);
  g29604 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output17(1), B1 => n_602, B2 => snake_output21(1), ZN => n_713);
  g29605 : AOI22D0BWP7T port map(A1 => n_617, A2 => snake_output8(1), B1 => n_512, B2 => snake_output9(1), ZN => n_712);
  g29606 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output18(2), B1 => n_502, B2 => snake_output20(2), ZN => n_711);
  g29607 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output17(2), B1 => n_602, B2 => snake_output21(2), ZN => n_710);
  g29608 : AOI22D0BWP7T port map(A1 => n_617, A2 => snake_output8(2), B1 => n_512, B2 => snake_output9(2), ZN => n_709);
  g29609 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output18(3), B1 => n_502, B2 => snake_output20(3), ZN => n_708);
  g29610 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output17(3), B1 => n_602, B2 => snake_output21(3), ZN => n_707);
  g29611 : AOI22D0BWP7T port map(A1 => n_617, A2 => snake_output8(3), B1 => n_512, B2 => snake_output9(3), ZN => n_706);
  g29612 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output18(4), B1 => n_502, B2 => snake_output20(4), ZN => n_705);
  g29613 : AOI22D0BWP7T port map(A1 => n_596, A2 => snake_output17(4), B1 => n_602, B2 => snake_output21(4), ZN => n_704);
  g29614 : AOI22D0BWP7T port map(A1 => n_617, A2 => snake_output8(4), B1 => n_512, B2 => snake_output9(4), ZN => n_703);
  g29615 : ND2D0BWP7T port map(A1 => n_699, A2 => n_1740, ZN => n_755);
  g29616 : NR3D0BWP7T port map(A1 => n_610, A2 => n_1699, A3 => n_156, ZN => n_754);
  g29619 : NR2D0BWP7T port map(A1 => n_193, A2 => n_684, ZN => n_752);
  g29620 : NR2D0BWP7T port map(A1 => n_193, A2 => n_686, ZN => n_751);
  g29621 : OAI21D0BWP7T port map(A1 => n_610, A2 => n_434, B => n_195, ZN => n_811);
  g29622 : AN2D1BWP7T port map(A1 => n_699, A2 => n_231, Z => n_750);
  g29626 : AN2D1BWP7T port map(A1 => n_699, A2 => n_227, Z => n_749);
  g29631 : OAI21D0BWP7T port map(A1 => n_610, A2 => n_1581, B => n_195, ZN => n_812);
  g29632 : CKND1BWP7T port map(I => n_700, ZN => n_701);
  g29633 : INVD0BWP7T port map(I => n_687, ZN => n_686);
  g29634 : CKND1BWP7T port map(I => n_685, ZN => n_684);
  g29635 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(2), B1 => n_539, B2 => snake_output3(2), ZN => n_683);
  g29636 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(1), B1 => n_539, B2 => snake_output3(1), ZN => n_682);
  g29637 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(0), B1 => n_539, B2 => snake_output3(0), ZN => n_681);
  g29638 : AOI22D0BWP7T port map(A1 => n_561, A2 => snake_output6(0), B1 => n_557, B2 => snake_output11(0), ZN => n_680);
  g29639 : AOI31D0BWP7T port map(A1 => n_1734, A2 => n_532, A3 => snake_output8(5), B => n_547, ZN => n_679);
  g29640 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(0), B1 => n_462, B2 => snake_output21(0), ZN => n_678);
  g29641 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(3), B1 => n_539, B2 => snake_output3(3), ZN => n_677);
  g29642 : ND4D0BWP7T port map(A1 => n_254, A2 => n_493, A3 => n_232, A4 => n_237, ZN => n_676);
  g29643 : AOI22D0BWP7T port map(A1 => n_540, A2 => snake_output4(4), B1 => n_539, B2 => snake_output3(4), ZN => n_675);
  g29644 : NR2D0BWP7T port map(A1 => n_610, A2 => n_438, ZN => n_700);
  g29645 : NR2D0BWP7T port map(A1 => n_619, A2 => corner_count(1), ZN => n_699);
  g29647 : INR2D0BWP7T port map(A1 => n_622, B1 => n_193, ZN => n_698);
  g29648 : NR2D0BWP7T port map(A1 => n_193, A2 => n_601, ZN => n_697);
  g29649 : NR3D0BWP7T port map(A1 => n_193, A2 => n_477, A3 => n_544, ZN => n_696);
  g29650 : NR2D0BWP7T port map(A1 => n_193, A2 => n_595, ZN => n_695);
  g29651 : NR2D0BWP7T port map(A1 => n_619, A2 => n_429, ZN => n_694);
  g29654 : NR2D0BWP7T port map(A1 => n_619, A2 => n_430, ZN => n_693);
  g29659 : OAI21D0BWP7T port map(A1 => n_541, A2 => n_217, B => n_195, ZN => n_765);
  g29660 : OAI21D0BWP7T port map(A1 => n_541, A2 => n_220, B => n_195, ZN => n_763);
  g29661 : AOI21D0BWP7T port map(A1 => n_565, A2 => n_212, B => n_194, ZN => n_762);
  g29662 : AOI21D0BWP7T port map(A1 => n_565, A2 => n_222, B => n_194, ZN => n_761);
  g29663 : AOI21D0BWP7T port map(A1 => n_564, A2 => n_222, B => n_194, ZN => n_759);
  g29665 : OAI21D0BWP7T port map(A1 => n_541, A2 => n_211, B => n_195, ZN => n_764);
  g29667 : IAO21D0BWP7T port map(A1 => n_566, A2 => n_220, B => n_194, ZN => n_757);
  g29669 : OAI21D0BWP7T port map(A1 => n_563, A2 => n_217, B => n_195, ZN => n_756);
  g29670 : AOI21D0BWP7T port map(A1 => n_565, A2 => n_218, B => n_194, ZN => n_758);
  g29672 : OAI21D0BWP7T port map(A1 => n_563, A2 => n_220, B => n_195, ZN => n_702);
  g29673 : AOI21D0BWP7T port map(A1 => n_564, A2 => n_212, B => n_194, ZN => n_760);
  g29674 : IOA21D0BWP7T port map(A1 => n_542, A2 => n_222, B => n_195, ZN => n_766);
  g29676 : NR2D0BWP7T port map(A1 => n_623, A2 => corner_count(0), ZN => n_692);
  g29677 : NR2D0BWP7T port map(A1 => n_623, A2 => n_146, ZN => n_691);
  g29678 : INR2D0BWP7T port map(A1 => n_425, B1 => n_619, ZN => n_690);
  g29679 : NR2D0BWP7T port map(A1 => n_619, A2 => n_428, ZN => n_689);
  g29680 : INR2D0BWP7T port map(A1 => n_622, B1 => n_478, ZN => n_688);
  g29681 : AN3D0BWP7T port map(A1 => n_477, A2 => n_544, A3 => n_420, Z => n_687);
  g29682 : NR3D0BWP7T port map(A1 => n_524, A2 => n_478, A3 => n_545, ZN => n_685);
  g29683 : AOI22D0BWP7T port map(A1 => n_546, A2 => snake_output17(5), B1 => n_462, B2 => snake_output22(5), ZN => n_672);
  g29684 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(0), B1 => n_496, B2 => snake_output1(0), ZN => n_671);
  g29685 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output11(0), B1 => n_418, B2 => snake_output14(0), ZN => n_670);
  g29686 : AOI22D0BWP7T port map(A1 => n_514, A2 => snake_output12(0), B1 => n_550, B2 => snake_output13(0), ZN => n_669);
  g29687 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(0), B1 => n_462, B2 => snake_output20(0), ZN => n_668);
  g29688 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output10(0), B1 => n_514, B2 => snake_output11(0), ZN => n_667);
  g29689 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(1), B1 => n_462, B2 => snake_output21(1), ZN => n_666);
  g29690 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output23(1), B1 => n_559, B2 => snake_output16(1), ZN => n_665);
  g29691 : AOI22D0BWP7T port map(A1 => n_543, A2 => snake_output24(5), B1 => n_475, B2 => snake_output16(5), ZN => n_664);
  g29692 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(1), B1 => n_496, B2 => snake_output1(1), ZN => n_663);
  g29693 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output14(5), B1 => n_418, B2 => snake_output15(5), ZN => n_662);
  g29694 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output11(1), B1 => n_418, B2 => snake_output14(1), ZN => n_661);
  g29695 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output12(5), B1 => n_514, B2 => snake_output13(5), ZN => n_660);
  g29696 : AOI22D0BWP7T port map(A1 => n_514, A2 => snake_output12(1), B1 => n_550, B2 => snake_output13(1), ZN => n_659);
  g29697 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(1), B1 => n_462, B2 => snake_output20(1), ZN => n_658);
  g29698 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output10(1), B1 => n_514, B2 => snake_output11(1), ZN => n_657);
  g29699 : AOI22D0BWP7T port map(A1 => n_510, A2 => snake_output1(1), B1 => n_532, B2 => snake_output5(1), ZN => n_656);
  g29700 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(2), B1 => n_462, B2 => snake_output21(2), ZN => n_655);
  g29701 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output23(2), B1 => n_559, B2 => snake_output16(2), ZN => n_654);
  g29702 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(2), B1 => n_496, B2 => snake_output1(2), ZN => n_653);
  g29703 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output1(5), B1 => n_507, B2 => snake_output0(5), ZN => n_652);
  g29704 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output11(2), B1 => n_418, B2 => snake_output14(2), ZN => n_651);
  g29705 : AOI22D0BWP7T port map(A1 => n_514, A2 => snake_output12(2), B1 => n_550, B2 => snake_output13(2), ZN => n_650);
  g29706 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(2), B1 => n_462, B2 => snake_output20(2), ZN => n_649);
  g29707 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output12(2), B1 => n_418, B2 => snake_output13(2), ZN => n_648);
  g29708 : AOI22D0BWP7T port map(A1 => n_510, A2 => snake_output1(2), B1 => n_532, B2 => snake_output5(2), ZN => n_647);
  g29709 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(3), B1 => n_462, B2 => snake_output21(3), ZN => n_646);
  g29710 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output23(3), B1 => n_559, B2 => snake_output16(3), ZN => n_645);
  g29711 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(3), B1 => n_496, B2 => snake_output1(3), ZN => n_644);
  g29712 : AOI22D0BWP7T port map(A1 => n_514, A2 => snake_output12(3), B1 => n_550, B2 => snake_output13(3), ZN => n_643);
  g29713 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(3), B1 => n_462, B2 => snake_output20(3), ZN => n_642);
  g29714 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output12(3), B1 => n_418, B2 => snake_output13(3), ZN => n_641);
  g29715 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output4(3), B1 => n_532, B2 => snake_output5(3), ZN => n_640);
  g29716 : AOI22D0BWP7T port map(A1 => n_534, A2 => snake_output19(4), B1 => n_462, B2 => snake_output21(4), ZN => n_639);
  g29717 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output23(4), B1 => n_559, B2 => snake_output16(4), ZN => n_638);
  g29718 : AOI22D0BWP7T port map(A1 => n_555, A2 => snake_output0(4), B1 => n_496, B2 => snake_output1(4), ZN => n_637);
  g29719 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output11(4), B1 => n_418, B2 => snake_output14(4), ZN => n_636);
  g29720 : AOI22D0BWP7T port map(A1 => n_514, A2 => snake_output12(4), B1 => n_550, B2 => snake_output13(4), ZN => n_635);
  g29721 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output22(4), B1 => n_462, B2 => snake_output20(4), ZN => n_634);
  g29722 : AOI22D0BWP7T port map(A1 => n_550, A2 => snake_output12(4), B1 => n_418, B2 => snake_output13(4), ZN => n_633);
  g29723 : AOI22D0BWP7T port map(A1 => n_552, A2 => snake_output11(3), B1 => n_418, B2 => snake_output14(3), ZN => n_632);
  g29724 : AOI22D0BWP7T port map(A1 => n_510, A2 => snake_output1(4), B1 => n_532, B2 => snake_output5(4), ZN => n_631);
  g29725 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output6(5), B1 => n_532, B2 => snake_output7(5), ZN => n_630);
  g29726 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(0), B1 => n_550, B2 => snake_output12(0), ZN => n_629);
  g29727 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(1), B1 => n_550, B2 => snake_output12(1), ZN => n_628);
  g29728 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(2), B1 => n_552, B2 => snake_output10(2), ZN => n_627);
  g29729 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(3), B1 => n_552, B2 => snake_output10(3), ZN => n_626);
  g29730 : AOI22D0BWP7T port map(A1 => n_503, A2 => snake_output15(4), B1 => n_552, B2 => snake_output10(4), ZN => n_625);
  g29731 : AOI22D0BWP7T port map(A1 => n_553, A2 => snake_output23(0), B1 => n_559, B2 => snake_output16(0), ZN => n_624);
  g29733 : CKND1BWP7T port map(I => n_602, ZN => n_601);
  g29734 : OAI31D0BWP7T port map(A1 => N(0), A2 => n_230, A3 => n_423, B => n_232, ZN => n_600);
  g29735 : AOI31D0BWP7T port map(A1 => n_485, A2 => N(0), A3 => snake_output1(5), B => n_489, ZN => n_599);
  g29736 : ND2D0BWP7T port map(A1 => n_536, A2 => n_228, ZN => n_623);
  g29737 : NR2D0BWP7T port map(A1 => n_523, A2 => n_545, ZN => n_622);
  g29738 : AN2D1BWP7T port map(A1 => n_478, A2 => n_545, Z => n_621);
  g29739 : INR2D0BWP7T port map(A1 => n_546, B1 => n_193, ZN => n_620);
  g29740 : ND2D0BWP7T port map(A1 => n_535, A2 => n_463, ZN => n_619);
  g29741 : INR2D0BWP7T port map(A1 => n_554, B1 => n_193, ZN => n_618);
  g29742 : INR2D0BWP7T port map(A1 => n_554, B1 => n_478, ZN => n_617);
  g29743 : NR2D0BWP7T port map(A1 => n_193, A2 => n_549, ZN => n_616);
  g29744 : NR2D0BWP7T port map(A1 => n_193, A2 => n_531, ZN => n_615);
  g29745 : INR2D0BWP7T port map(A1 => n_555, B1 => n_193, ZN => n_614);
  g29746 : NR2D0BWP7T port map(A1 => n_193, A2 => n_551, ZN => n_613);
  g29747 : NR2D0BWP7T port map(A1 => n_193, A2 => n_533, ZN => n_612);
  g29748 : AOI211D0BWP7T port map(A1 => n_485, A2 => N(4), B => n_464, C => n_508, ZN => n_611);
  g29750 : ND2D0BWP7T port map(A1 => n_529, A2 => n_1698, ZN => n_610);
  g29751 : INR2D0BWP7T port map(A1 => n_425, B1 => n_535, ZN => n_609);
  g29753 : NR2D0BWP7T port map(A1 => n_535, A2 => n_428, ZN => n_608);
  g29755 : NR2D0BWP7T port map(A1 => n_535, A2 => n_435, ZN => n_607);
  g29758 : NR2D0BWP7T port map(A1 => n_535, A2 => n_436, ZN => n_606);
  g29759 : NR2D0BWP7T port map(A1 => n_535, A2 => n_430, ZN => n_605);
  g29760 : NR2D0BWP7T port map(A1 => n_535, A2 => n_463, ZN => n_604);
  g29762 : NR3D0BWP7T port map(A1 => n_429, A2 => n_536, A3 => n_463, ZN => n_603);
  g29763 : OAI21D0BWP7T port map(A1 => n_522, A2 => n_1700, B => n_195, ZN => n_674);
  g29764 : NR4D1BWP7T port map(A1 => n_477, A2 => n_466, A3 => n_421, A4 => N(0), ZN => n_602);
  g29765 : INVD0BWP7T port map(I => n_596, ZN => n_595);
  g29766 : AOI22D0BWP7T port map(A1 => n_498, A2 => snake_output2(3), B1 => n_510, B2 => snake_output1(3), ZN => n_594);
  g29767 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(1), B1 => n_519, B2 => snake_output11(1), ZN => n_593);
  g29768 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(1), B1 => n_505, B2 => snake_output13(1), ZN => n_592);
  g29769 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(2), B1 => n_519, B2 => snake_output11(2), ZN => n_591);
  g29770 : AOI22D0BWP7T port map(A1 => n_512, A2 => snake_output10(0), B1 => n_475, B2 => snake_output15(0), ZN => n_590);
  g29771 : AOI22D0BWP7T port map(A1 => n_506, A2 => snake_output16(0), B1 => n_502, B2 => snake_output19(0), ZN => n_589);
  g29772 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output4(0), B1 => n_496, B2 => snake_output0(0), ZN => n_588);
  g29773 : AOI22D0BWP7T port map(A1 => n_512, A2 => snake_output10(1), B1 => n_475, B2 => snake_output15(1), ZN => n_587);
  g29774 : AOI22D0BWP7T port map(A1 => n_506, A2 => snake_output16(1), B1 => n_502, B2 => snake_output19(1), ZN => n_586);
  g29775 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output4(1), B1 => n_496, B2 => snake_output0(1), ZN => n_585);
  g29776 : AOI22D0BWP7T port map(A1 => n_498, A2 => n_1167, B1 => n_510, B2 => snake_output3(5), ZN => n_584);
  g29777 : AOI22D0BWP7T port map(A1 => n_512, A2 => snake_output10(2), B1 => n_475, B2 => snake_output15(2), ZN => n_583);
  g29778 : AOI22D0BWP7T port map(A1 => n_506, A2 => snake_output16(2), B1 => n_502, B2 => snake_output19(2), ZN => n_582);
  g29779 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output4(2), B1 => n_496, B2 => snake_output0(2), ZN => n_581);
  g29780 : AOI22D0BWP7T port map(A1 => n_512, A2 => snake_output10(3), B1 => n_475, B2 => snake_output15(3), ZN => n_580);
  g29781 : AOI22D0BWP7T port map(A1 => n_506, A2 => snake_output16(3), B1 => n_502, B2 => snake_output19(3), ZN => n_579);
  g29782 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(2), B1 => n_505, B2 => snake_output13(2), ZN => n_578);
  g29783 : AOI22D0BWP7T port map(A1 => n_512, A2 => snake_output10(4), B1 => n_475, B2 => snake_output15(4), ZN => n_577);
  g29784 : AOI22D0BWP7T port map(A1 => n_506, A2 => snake_output16(4), B1 => n_502, B2 => snake_output19(4), ZN => n_576);
  g29785 : AOI22D0BWP7T port map(A1 => n_500, A2 => snake_output4(4), B1 => n_496, B2 => snake_output0(4), ZN => n_575);
  g29786 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(5), B1 => n_519, B2 => snake_output11(5), ZN => n_574);
  g29787 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(5), B1 => n_505, B2 => snake_output13(5), ZN => n_573);
  g29788 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(4), B1 => n_505, B2 => snake_output13(4), ZN => n_572);
  g29789 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(4), B1 => n_519, B2 => snake_output11(4), ZN => n_571);
  g29790 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(3), B1 => n_505, B2 => snake_output13(3), ZN => n_570);
  g29791 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(3), B1 => n_519, B2 => snake_output11(3), ZN => n_569);
  g29792 : AOI22D0BWP7T port map(A1 => n_504, A2 => snake_output10(0), B1 => n_519, B2 => snake_output11(0), ZN => n_568);
  g29793 : AOI22D0BWP7T port map(A1 => n_520, A2 => snake_output12(0), B1 => n_505, B2 => snake_output13(0), ZN => n_567);
  g29794 : AO21D0BWP7T port map(A1 => n_192, A2 => n_507, B => n_1737, Z => n_597);
  g29795 : IAO21D0BWP7T port map(A1 => n_522, A2 => n_150, B => n_194, ZN => n_673);
  g29797 : INR4D1BWP7T port map(A1 => n_466, B1 => N(0), B2 => n_421, B3 => n_477, ZN => n_596);
  g29798 : CKND1BWP7T port map(I => n_565, ZN => n_566);
  g29799 : CKND1BWP7T port map(I => n_564, ZN => n_563);
  g29800 : CKND1BWP7T port map(I => n_552, ZN => n_551);
  g29801 : CKND1BWP7T port map(I => n_550, ZN => n_549);
  g29803 : NR2D0BWP7T port map(A1 => n_492, A2 => n_230, ZN => n_547);
  g29804 : NR2D0BWP7T port map(A1 => n_525, A2 => n_1701, ZN => n_565);
  g29805 : NR2D0BWP7T port map(A1 => n_525, A2 => n_156, ZN => n_564);
  g29806 : NR2D0BWP7T port map(A1 => n_523, A2 => n_479, ZN => n_562);
  g29807 : NR2D0BWP7T port map(A1 => n_193, A2 => n_499, ZN => n_561);
  g29808 : NR2D0BWP7T port map(A1 => n_193, A2 => n_501, ZN => n_560);
  g29809 : AN2D1BWP7T port map(A1 => n_503, A2 => N(4), Z => n_559);
  g29810 : NR2D0BWP7T port map(A1 => n_193, A2 => n_513, ZN => n_558);
  g29811 : NR2D0BWP7T port map(A1 => n_193, A2 => n_511, ZN => n_557);
  g29812 : INR2D0BWP7T port map(A1 => n_515, B1 => n_193, ZN => n_556);
  g29813 : AN2D1BWP7T port map(A1 => n_503, A2 => n_477, Z => n_555);
  g29814 : NR2D0BWP7T port map(A1 => n_521, A2 => n_224, ZN => n_554);
  g29815 : NR2D0BWP7T port map(A1 => n_524, A2 => n_479, ZN => n_553);
  g29816 : INR2XD0BWP7T port map(A1 => n_226, B1 => n_521, ZN => n_552);
  g29817 : NR2D1BWP7T port map(A1 => n_521, A2 => n_221, ZN => n_550);
  g29818 : INVD0BWP7T port map(I => n_544, ZN => n_543);
  g29819 : CKND1BWP7T port map(I => n_541, ZN => n_542);
  g29820 : INVD1BWP7T port map(I => n_536, ZN => n_535);
  g29821 : CKND1BWP7T port map(I => n_534, ZN => n_533);
  g29822 : INVD1BWP7T port map(I => n_531, ZN => n_532);
  g29823 : INR4D0BWP7T port map(A1 => n_452, B1 => n_1734, B2 => n_1739, B3 => n_1737, ZN => n_530);
  g29824 : NR4D0BWP7T port map(A1 => n_469, A2 => n_1695, A3 => n_1696, A4 => n_1697, ZN => n_529);
  g29825 : INR4D0BWP7T port map(A1 => n_449, B1 => corner_count(31), B2 => corner_count(30), B3 => corner_count(29), ZN => n_528);
  g29826 : AOI22D0BWP7T port map(A1 => n_475, A2 => snake_output14(0), B1 => n_418, B2 => snake_output13(0), ZN => n_527);
  g29827 : AOI31D0BWP7T port map(A1 => n_214, A2 => N(3), A3 => snake_output24(5), B => n_491, ZN => n_526);
  g29828 : AN3D0BWP7T port map(A1 => n_476, A2 => n_468, A3 => n_466, Z => n_546);
  g29829 : OAI21D0BWP7T port map(A1 => n_484, A2 => n_149, B => n_424, ZN => n_545);
  g29830 : AOI21D0BWP7T port map(A1 => n_488, A2 => N(3), B => n_418, ZN => n_544);
  g29831 : IND3D0BWP7T port map(A1 => n_1699, B1 => n_1701, B2 => n_481, ZN => n_541);
  g29832 : NR2D0BWP7T port map(A1 => n_193, A2 => n_497, ZN => n_540);
  g29833 : NR2D0BWP7T port map(A1 => n_193, A2 => n_509, ZN => n_539);
  g29834 : NR3D0BWP7T port map(A1 => n_193, A2 => n_474, A3 => n_477, ZN => n_538);
  g29835 : NR2D0BWP7T port map(A1 => n_193, A2 => n_495, ZN => n_537);
  g29836 : IAO21D0BWP7T port map(A1 => n_482, A2 => n_434, B => n_194, ZN => n_598);
  g29837 : CKXOR2D0BWP7T port map(A1 => corner_count(4), A2 => n_419, Z => n_536);
  g29838 : NR3D0BWP7T port map(A1 => n_467, A2 => n_466, A3 => n_147, ZN => n_534);
  g29839 : ND3D0BWP7T port map(A1 => n_426, A2 => n_147, A3 => N(3), ZN => n_531);
  g29840 : CKND1BWP7T port map(I => n_514, ZN => n_513);
  g29841 : CKND1BWP7T port map(I => n_512, ZN => n_511);
  g29842 : CKND1BWP7T port map(I => n_510, ZN => n_509);
  g29843 : NR2D0BWP7T port map(A1 => n_485, A2 => N(4), ZN => n_508);
  g29844 : ND2D0BWP7T port map(A1 => n_481, A2 => n_1699, ZN => n_525);
  g29845 : OR2D0BWP7T port map(A1 => n_467, A2 => n_486, Z => n_524);
  g29846 : ND2D0BWP7T port map(A1 => n_468, A2 => n_487, ZN => n_523);
  g29847 : IND2D0BWP7T port map(A1 => n_438, B1 => n_481, ZN => n_522);
  g29848 : IND2D0BWP7T port map(A1 => n_464, B1 => N(0), ZN => n_521);
  g29849 : INR2D0BWP7T port map(A1 => n_425, B1 => n_463, ZN => n_520);
  g29850 : NR2D0BWP7T port map(A1 => n_435, A2 => n_463, ZN => n_519);
  g29851 : INR2D0BWP7T port map(A1 => n_419, B1 => n_146, ZN => n_518);
  g29852 : INR2D0BWP7T port map(A1 => n_419, B1 => corner_count(0), ZN => n_517);
  g29853 : NR2D0BWP7T port map(A1 => n_428, A2 => n_463, ZN => n_516);
  g29854 : NR2D0BWP7T port map(A1 => n_487, A2 => n_439, ZN => n_515);
  g29855 : INR2XD0BWP7T port map(A1 => n_420, B1 => n_464, ZN => n_514);
  g29856 : NR2D1BWP7T port map(A1 => n_464, A2 => n_433, ZN => n_512);
  g29857 : NR2D1BWP7T port map(A1 => n_478, A2 => n_437, ZN => n_510);
  g29858 : INVD1BWP7T port map(I => n_501, ZN => n_502);
  g29859 : CKND1BWP7T port map(I => n_500, ZN => n_499);
  g29860 : CKND1BWP7T port map(I => n_498, ZN => n_497);
  g29861 : CKND1BWP7T port map(I => n_496, ZN => n_495);
  g29862 : AOI33D0BWP7T port map(A1 => n_432, A2 => n_214, A3 => snake_output20(5), B1 => n_420, B2 => n_223, B3 => snake_output14(5), ZN => n_494);
  g29863 : MAOI22D0BWP7T port map(A1 => n_1572, A2 => n_448, B1 => n_154, B2 => send_corner_flag, ZN => n_493);
  g29864 : AOI31D0BWP7T port map(A1 => n_420, A2 => n_149, A3 => snake_output6(5), B => n_457, ZN => n_492);
  g29865 : NR3D0BWP7T port map(A1 => n_460, A2 => n_224, A3 => N(0), ZN => n_491);
  g29866 : AOI22D0BWP7T port map(A1 => n_442, A2 => n_427, B1 => n_458, B2 => snake_output12(5), ZN => n_490);
  g29867 : OAI32D0BWP7T port map(A1 => n_153, A2 => n_215, A3 => n_239, B1 => n_144, B2 => n_437, ZN => n_489);
  g29868 : NR2D0BWP7T port map(A1 => n_474, A2 => n_476, ZN => n_507);
  g29869 : NR2D0BWP7T port map(A1 => n_479, A2 => n_441, ZN => n_506);
  g29870 : NR2D0BWP7T port map(A1 => n_430, A2 => n_463, ZN => n_505);
  g29871 : NR2D0BWP7T port map(A1 => n_436, A2 => n_463, ZN => n_504);
  g29872 : AN3D0BWP7T port map(A1 => n_464, A2 => n_468, A3 => n_221, Z => n_503);
  g29873 : ND2D0BWP7T port map(A1 => n_476, A2 => n_420, ZN => n_501);
  g29874 : NR3D0BWP7T port map(A1 => n_478, A2 => n_421, A3 => n_431, ZN => n_500);
  g29875 : NR3D0BWP7T port map(A1 => n_476, A2 => n_422, A3 => n_431, ZN => n_498);
  g29876 : NR2D1BWP7T port map(A1 => n_478, A2 => n_441, ZN => n_496);
  g29877 : CKND1BWP7T port map(I => n_426, ZN => n_488);
  g29879 : INVD0BWP7T port map(I => n_486, ZN => n_487);
  g29880 : CKND1BWP7T port map(I => n_423, ZN => n_485);
  g29881 : HA1D0BWP7T port map(A => n_148, B => n_210, CO => n_484, S => n_486);
  g29902 : CKND1BWP7T port map(I => n_481, ZN => n_482);
  g29903 : INVD1BWP7T port map(I => n_479, ZN => n_478);
  g29904 : INVD1BWP7T port map(I => n_477, ZN => n_476);
  g29905 : CKND1BWP7T port map(I => n_475, ZN => n_474);
  g29913 : AOI22D0BWP7T port map(A1 => n_418, A2 => snake_output16(5), B1 => n_420, B2 => snake_output22(5), ZN => n_473);
  g29918 : MAOI22D0BWP7T port map(A1 => n_427, A2 => snake_output15(5), B1 => n_440, B2 => n_145, ZN => n_472);
  g29920 : AOI222D0BWP7T port map(A1 => n_219, A2 => snake_output17(5), B1 => n_226, B2 => snake_output21(5), C1 => n_225, C2 => snake_output19(5), ZN => n_471);
  g29921 : NR2D0BWP7T port map(A1 => n_469, A2 => n_1582, ZN => n_481);
  g29922 : NR2D0BWP7T port map(A1 => n_193, A2 => n_461, ZN => n_480);
  g29923 : MAOI22D0BWP7T port map(A1 => n_424, A2 => N(4), B1 => n_424, B2 => N(4), ZN => n_479);
  g29925 : AOI22D0BWP7T port map(A1 => n_418, A2 => n_147, B1 => n_417, B2 => N(4), ZN => n_477);
  g29926 : NR2D1BWP7T port map(A1 => n_467, A2 => n_215, ZN => n_475);
  g29956 : CKND1BWP7T port map(I => n_462, ZN => n_461);
  g29957 : AOI22D0BWP7T port map(A1 => n_214, A2 => snake_output18(5), B1 => n_223, B2 => snake_output10(5), ZN => n_460);
  g29958 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(4), B1 => n_207, B2 => snake_output0(4), ZN => n_459);
  g29959 : INR2D0BWP7T port map(A1 => n_223, B1 => n_433, ZN => n_458);
  g29960 : NR2D0BWP7T port map(A1 => n_431, A2 => n_238, ZN => n_457);
  g29961 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(3), B1 => n_207, B2 => snake_output0(3), ZN => n_456);
  g29962 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(1), B1 => n_207, B2 => snake_output0(1), ZN => n_455);
  g29963 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(0), B1 => n_207, B2 => snake_output0(0), ZN => n_454);
  g29964 : AOI22D0BWP7T port map(A1 => n_209, A2 => head(2), B1 => n_1737, B2 => head(7), ZN => n_453);
  g29965 : NR4D0BWP7T port map(A1 => n_1579, A2 => n_1735, A3 => n_1736, A4 => n_1738, ZN => n_452);
  g29966 : AO221D0BWP7T port map(A1 => n_1703, A2 => n_146, B1 => FE_OFN3_n_1704, B2 => new_corner_count(0), C => n_1739, Z => n_451);
  g29967 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(4), B1 => n_207, B2 => head(9), ZN => n_450);
  g29968 : NR4D0BWP7T port map(A1 => corner_count(16), A2 => corner_count(15), A3 => corner_count(14), A4 => corner_count(13), ZN => n_449);
  g29969 : AO211D0BWP7T port map(A1 => n_1273, A2 => n_1742, B => n_1575, C => new_head_flag, Z => n_448);
  g29970 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(3), B1 => n_207, B2 => head(8), ZN => n_447);
  g29971 : IIND4D0BWP7T port map(A1 => n_1573, A2 => n_1574, B1 => n_1572, B2 => n_1585, ZN => n_446);
  g29972 : AOI22D0BWP7T port map(A1 => n_207, A2 => head(7), B1 => n_1737, B2 => head(2), ZN => n_445);
  g29973 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(1), B1 => n_207, B2 => head(6), ZN => n_444);
  g29974 : AOI22D0BWP7T port map(A1 => n_209, A2 => snake_output0(0), B1 => n_207, B2 => head(5), ZN => n_443);
  g29975 : AO22D0BWP7T port map(A1 => n_219, A2 => snake_output9(5), B1 => snake_output11(5), B2 => n_225, Z => n_442);
  g29976 : OAI211D0BWP7T port map(A1 => n_1670, A2 => n_1703, B => n_1580, C => n_187, ZN => n_469);
  g29978 : NR2D0BWP7T port map(A1 => n_422, A2 => N(0), ZN => n_468);
  g29979 : ND2D0BWP7T port map(A1 => n_421, A2 => N(0), ZN => n_467);
  g29981 : AOI21D0BWP7T port map(A1 => n_216, A2 => N(2), B => n_426, ZN => n_466);
  g29982 : NR2D0BWP7T port map(A1 => n_193, A2 => n_417, ZN => n_465);
  g29983 : OA21D0BWP7T port map(A1 => n_219, A2 => n_149, B => n_423, Z => n_464);
  g29984 : AOI21D0BWP7T port map(A1 => n_229, A2 => corner_count(3), B => n_419, ZN => n_463);
  g29985 : NR2D1BWP7T port map(A1 => n_439, A2 => n_148, ZN => n_462);
  g29986 : NR4D0BWP7T port map(A1 => n_1739, A2 => n_1734, A3 => n_1662, A4 => n_1736, ZN => n_483);
  g29987 : INVD0BWP7T port map(I => n_433, ZN => n_432);
  g29988 : INVD1BWP7T port map(I => n_422, ZN => n_421);
  g29989 : INVD1BWP7T port map(I => n_418, ZN => n_417);
  g29995 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift9(1), B => n_201, ZN => n_416);
  g29996 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift8(5), B => n_197, ZN => n_415);
  g29997 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift8(3), B => n_198, ZN => n_414);
  g29998 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift5(3), B => n_198, ZN => n_413);
  g29999 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift8(1), B => n_201, ZN => n_412);
  g30000 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift7(5), B => n_197, ZN => n_411);
  g30001 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(5), B => n_197, ZN => n_410);
  g30002 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift7(4), B => n_196, ZN => n_409);
  g30003 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift7(3), B => n_198, ZN => n_408);
  g30004 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift16(0), B => n_199, ZN => n_407);
  g30005 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift6(0), B => n_199, ZN => n_406);
  g30006 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift7(1), B => n_201, ZN => n_405);
  g30007 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift6(4), B => n_196, ZN => n_404);
  g30008 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift6(3), B => n_198, ZN => n_403);
  g30009 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift6(2), B => n_200, ZN => n_402);
  g30010 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift4(1), B => n_201, ZN => n_401);
  g30011 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift8(2), B => n_200, ZN => n_400);
  g30012 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift6(1), B => n_201, ZN => n_399);
  g30013 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift4(2), B => n_200, ZN => n_398);
  g30014 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift8(0), B => n_199, ZN => n_397);
  g30015 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift2(0), B => n_199, ZN => n_396);
  g30016 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift4(4), B => n_196, ZN => n_395);
  g30017 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift4(0), B => n_199, ZN => n_394);
  g30018 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(1), B => n_201, ZN => n_393);
  g30019 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift19(0), B => n_199, ZN => n_392);
  g30020 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift19(1), B => n_201, ZN => n_391);
  g30021 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift19(2), B => n_200, ZN => n_390);
  g30022 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift19(3), B => n_198, ZN => n_389);
  g30023 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(2), B => n_200, ZN => n_388);
  g30024 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift19(4), B => n_196, ZN => n_387);
  g30025 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(3), B => n_198, ZN => n_386);
  g30026 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift19(5), B => n_197, ZN => n_385);
  g30027 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift20(0), B => n_199, ZN => n_384);
  g30028 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift20(1), B => n_201, ZN => n_383);
  g30029 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift20(2), B => n_200, ZN => n_382);
  g30030 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(4), B => n_196, ZN => n_381);
  g30031 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift20(3), B => n_198, ZN => n_380);
  g30032 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift20(4), B => n_196, ZN => n_379);
  g30033 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift20(5), B => n_197, ZN => n_378);
  g30034 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift21(0), B => n_199, ZN => n_377);
  g30035 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(0), B => n_199, ZN => n_376);
  g30036 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift4(5), B => n_197, ZN => n_375);
  g30037 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(5), B => n_197, ZN => n_374);
  g30038 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift21(1), B => n_201, ZN => n_373);
  g30039 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift21(2), B => n_200, ZN => n_372);
  g30040 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift21(3), B => n_198, ZN => n_371);
  g30041 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(2), B => n_200, ZN => n_370);
  g30042 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift22(0), B => n_199, ZN => n_369);
  g30043 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift22(1), B => n_201, ZN => n_368);
  g30044 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(3), B => n_198, ZN => n_367);
  g30045 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift22(2), B => n_200, ZN => n_366);
  g30046 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift22(4), B => n_196, ZN => n_365);
  g30047 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift22(5), B => n_197, ZN => n_364);
  g30048 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(4), B => n_196, ZN => n_363);
  g30049 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift23(0), B => n_199, ZN => n_362);
  g30050 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift23(1), B => n_201, ZN => n_361);
  g30051 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift8(4), B => n_196, ZN => n_360);
  g30052 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift23(4), B => n_196, ZN => n_359);
  g30053 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift23(3), B => n_198, ZN => n_358);
  g30054 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift23(5), B => n_197, ZN => n_357);
  g30055 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift3(5), B => n_197, ZN => n_356);
  g30056 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift2(2), B => n_200, ZN => n_355);
  g30057 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift5(4), B => n_196, ZN => n_354);
  g30058 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(1), B => n_201, ZN => n_353);
  g30059 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(4), B => n_196, ZN => n_352);
  g30060 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift23(2), B => n_200, ZN => n_351);
  g30061 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift2(5), B => n_197, ZN => n_350);
  g30062 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift3(0), B => n_199, ZN => n_349);
  g30063 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift1(1), B => n_201, ZN => n_348);
  g30064 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift21(5), B => n_197, ZN => n_347);
  g30065 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift21(4), B => n_196, ZN => n_346);
  g30066 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift3(2), B => n_200, ZN => n_345);
  g30067 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(3), B => n_198, ZN => n_344);
  g30068 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(4), B => n_196, ZN => n_343);
  g30069 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift7(0), B => n_199, ZN => n_342);
  g30070 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift22(3), B => n_198, ZN => n_341);
  g30071 : OR2D0BWP7T port map(A1 => n_210, A2 => n_215, Z => n_441);
  g30072 : ND2D0BWP7T port map(A1 => n_214, A2 => N(0), ZN => n_440);
  g30073 : IND2D0BWP7T port map(A1 => n_210, B1 => N(4), ZN => n_439);
  g30074 : ND2D0BWP7T port map(A1 => n_235, A2 => n_146, ZN => n_438);
  g30075 : IND2D0BWP7T port map(A1 => n_216, B1 => n_234, ZN => n_437);
  g30076 : IND2D0BWP7T port map(A1 => corner_count(1), B1 => n_231, ZN => n_436);
  g30077 : IND2D0BWP7T port map(A1 => corner_count(1), B1 => n_227, ZN => n_435);
  g30078 : ND2D0BWP7T port map(A1 => n_235, A2 => n_218, ZN => n_434);
  g30079 : ND2D0BWP7T port map(A1 => n_226, A2 => n_152, ZN => n_433);
  g30080 : ND2D0BWP7T port map(A1 => n_234, A2 => N(0), ZN => n_431);
  g30081 : IND2D0BWP7T port map(A1 => n_233, B1 => corner_count(0), ZN => n_430);
  g30082 : ND2D0BWP7T port map(A1 => n_231, A2 => corner_count(1), ZN => n_429);
  g30083 : ND2D0BWP7T port map(A1 => n_227, A2 => corner_count(1), ZN => n_428);
  g30084 : AN2D1BWP7T port map(A1 => n_223, A2 => N(0), Z => n_427);
  g30085 : NR2D0BWP7T port map(A1 => n_216, A2 => N(2), ZN => n_426);
  g30086 : NR2D0BWP7T port map(A1 => n_233, A2 => corner_count(0), ZN => n_425);
  g30087 : IND2D0BWP7T port map(A1 => n_215, B1 => n_210, ZN => n_424);
  g30088 : ND2D0BWP7T port map(A1 => n_219, A2 => n_149, ZN => n_423);
  g30089 : ND2D0BWP7T port map(A1 => n_210, A2 => n_216, ZN => n_422);
  g30090 : NR2D0BWP7T port map(A1 => n_221, A2 => N(0), ZN => n_420);
  g30091 : NR2D0BWP7T port map(A1 => n_229, A2 => corner_count(3), ZN => n_419);
  g30092 : NR2D1BWP7T port map(A1 => n_215, A2 => n_216, ZN => n_418);
  g30093 : NR2XD1BWP7T port map(A1 => n_194, A2 => n_1703, ZN => n_470);
  g30094 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift9(2), B => n_200, ZN => n_340);
  g30095 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift9(3), B => n_198, ZN => n_339);
  g30096 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift9(4), B => n_196, ZN => n_338);
  g30097 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift9(5), B => n_197, ZN => n_337);
  g30098 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift10(0), B => n_199, ZN => n_336);
  g30099 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift4(3), B => n_198, ZN => n_335);
  g30100 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift10(1), B => n_201, ZN => n_334);
  g30101 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift10(2), B => n_200, ZN => n_333);
  g30102 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift10(3), B => n_198, ZN => n_332);
  g30103 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift10(4), B => n_196, ZN => n_331);
  g30104 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift10(5), B => n_197, ZN => n_330);
  g30105 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift11(0), B => n_199, ZN => n_329);
  g30106 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift9(0), B => n_199, ZN => n_328);
  g30107 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift11(1), B => n_201, ZN => n_327);
  g30108 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift11(2), B => n_200, ZN => n_326);
  g30109 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift11(3), B => n_198, ZN => n_325);
  g30110 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift11(4), B => n_196, ZN => n_324);
  g30111 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift11(5), B => n_197, ZN => n_323);
  g30112 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift12(0), B => n_199, ZN => n_322);
  g30113 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift5(0), B => n_199, ZN => n_321);
  g30114 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift12(1), B => n_201, ZN => n_320);
  g30115 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift7(2), B => n_200, ZN => n_319);
  g30116 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift12(2), B => n_200, ZN => n_318);
  g30117 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift12(3), B => n_198, ZN => n_317);
  g30118 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift12(4), B => n_196, ZN => n_316);
  g30119 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift12(5), B => n_197, ZN => n_315);
  g30120 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift13(0), B => n_199, ZN => n_314);
  g30121 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift13(1), B => n_201, ZN => n_313);
  g30122 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift13(2), B => n_200, ZN => n_312);
  g30123 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift13(3), B => n_198, ZN => n_311);
  g30124 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift13(4), B => n_196, ZN => n_310);
  g30125 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift13(5), B => n_197, ZN => n_309);
  g30126 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift6(5), B => n_197, ZN => n_308);
  g30127 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift14(0), B => n_199, ZN => n_307);
  g30128 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift14(1), B => n_201, ZN => n_306);
  g30129 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift14(2), B => n_200, ZN => n_305);
  g30130 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift14(3), B => n_198, ZN => n_304);
  g30131 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift14(4), B => n_196, ZN => n_303);
  g30132 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift14(5), B => n_197, ZN => n_302);
  g30133 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift15(0), B => n_199, ZN => n_301);
  g30134 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift15(1), B => n_201, ZN => n_300);
  g30135 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift15(2), B => n_200, ZN => n_299);
  g30136 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift3(1), B => n_201, ZN => n_298);
  g30137 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift15(3), B => n_198, ZN => n_297);
  g30138 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift15(4), B => n_196, ZN => n_296);
  g30139 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift15(5), B => n_197, ZN => n_295);
  g30140 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift2(3), B => n_198, ZN => n_294);
  g30141 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift16(1), B => n_201, ZN => n_293);
  g30142 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift16(2), B => n_200, ZN => n_292);
  g30143 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift16(3), B => n_198, ZN => n_291);
  g30144 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift16(4), B => n_196, ZN => n_290);
  g30145 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift16(5), B => n_197, ZN => n_289);
  g30146 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift5(5), B => n_197, ZN => n_288);
  g30147 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift17(0), B => n_199, ZN => n_287);
  g30148 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift5(2), B => n_200, ZN => n_286);
  g30149 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift17(1), B => n_201, ZN => n_285);
  g30150 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift5(1), B => n_201, ZN => n_284);
  g30151 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift17(2), B => n_200, ZN => n_283);
  g30152 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift17(3), B => n_198, ZN => n_282);
  g30153 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift17(4), B => n_196, ZN => n_281);
  g30154 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift17(5), B => n_197, ZN => n_280);
  g30155 : IOA21D0BWP7T port map(A1 => n_1704, A2 => shift0(0), B => n_199, ZN => n_279);
  g30156 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift18(0), B => n_199, ZN => n_278);
  g30157 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift18(1), B => n_201, ZN => n_277);
  g30158 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift18(2), B => n_200, ZN => n_276);
  g30159 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift18(3), B => n_198, ZN => n_275);
  g30160 : IOA21D0BWP7T port map(A1 => FE_OFN4_n_1704, A2 => shift18(4), B => n_196, ZN => n_274);
  g30161 : IOA21D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => shift18(5), B => n_197, ZN => n_273);
  g30162 : AO22D0BWP7T port map(A1 => n_1693, A2 => n_1703, B1 => new_corner_count(9), B2 => FE_OFN3_n_1704, Z => n_272);
  g30163 : AO22D0BWP7T port map(A1 => n_1692, A2 => n_1703, B1 => new_corner_count(10), B2 => FE_OFN3_n_1704, Z => n_271);
  g30164 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1698, B1 => new_corner_count(4), B2 => FE_OFN3_n_1704, Z => n_270);
  g30165 : MOAI22D0BWP7T port map(A1 => n_151, A2 => n_150, B1 => FE_OFN3_n_1704, B2 => new_corner_count(2), ZN => n_269);
  g30166 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1699, B1 => new_corner_count(3), B2 => FE_OFN3_n_1704, Z => n_268);
  g30167 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1697, B1 => new_corner_count(5), B2 => FE_OFN3_n_1704, Z => n_267);
  g30168 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1696, B1 => new_corner_count(6), B2 => FE_OFN3_n_1704, Z => n_266);
  g30169 : AO22D0BWP7T port map(A1 => n_1703, A2 => n_1695, B1 => new_corner_count(7), B2 => FE_OFN3_n_1704, Z => n_265);
  g30170 : AO22D0BWP7T port map(A1 => n_1694, A2 => n_1703, B1 => new_corner_count(8), B2 => FE_OFN3_n_1704, Z => n_264);
  g30171 : AO22D0BWP7T port map(A1 => n_1680, A2 => n_1703, B1 => new_corner_count(22), B2 => n_1704, Z => n_263);
  g30172 : AO22D0BWP7T port map(A1 => n_1691, A2 => n_1703, B1 => new_corner_count(11), B2 => FE_OFN3_n_1704, Z => n_262);
  g30173 : AO22D0BWP7T port map(A1 => n_1689, A2 => n_1703, B1 => new_corner_count(13), B2 => FE_OFN3_n_1704, Z => n_261);
  g30174 : AO22D0BWP7T port map(A1 => n_1684, A2 => n_1703, B1 => new_corner_count(18), B2 => FE_OFN3_n_1704, Z => n_260);
  g30175 : AO22D0BWP7T port map(A1 => n_1683, A2 => n_1703, B1 => new_corner_count(19), B2 => FE_OFN3_n_1704, Z => n_259);
  g30176 : AO22D0BWP7T port map(A1 => n_1679, A2 => n_1703, B1 => new_corner_count(23), B2 => n_1704, Z => n_258);
  g30177 : AO22D0BWP7T port map(A1 => n_1676, A2 => n_1703, B1 => new_corner_count(26), B2 => n_1704, Z => n_257);
  g30178 : AO22D0BWP7T port map(A1 => n_1675, A2 => n_1703, B1 => new_corner_count(27), B2 => n_1704, Z => n_256);
  g30179 : AO22D0BWP7T port map(A1 => n_1672, A2 => n_1703, B1 => new_corner_count(30), B2 => n_1704, Z => n_255);
  g30180 : NR4D0BWP7T port map(A1 => n_1731, A2 => n_1705, A3 => n_1718, A4 => n_1663, ZN => n_254);
  g30181 : AO22D0BWP7T port map(A1 => n_1685, A2 => n_1703, B1 => new_corner_count(17), B2 => FE_OFN3_n_1704, Z => n_253);
  g30182 : AO22D0BWP7T port map(A1 => n_1671, A2 => n_1703, B1 => new_corner_count(31), B2 => n_1704, Z => n_252);
  g30183 : MOAI22D0BWP7T port map(A1 => n_151, A2 => n_156, B1 => FE_OFN3_n_1704, B2 => new_corner_count(1), ZN => n_251);
  g30184 : AO22D0BWP7T port map(A1 => n_1690, A2 => n_1703, B1 => new_corner_count(12), B2 => FE_OFN3_n_1704, Z => n_250);
  g30185 : AO22D0BWP7T port map(A1 => n_1673, A2 => n_1703, B1 => new_corner_count(29), B2 => n_1704, Z => n_249);
  g30186 : AO22D0BWP7T port map(A1 => n_1681, A2 => n_1703, B1 => new_corner_count(21), B2 => FE_OFN3_n_1704, Z => n_248);
  g30187 : AO22D0BWP7T port map(A1 => n_1688, A2 => n_1703, B1 => new_corner_count(14), B2 => FE_OFN3_n_1704, Z => n_247);
  g30188 : AO22D0BWP7T port map(A1 => n_1674, A2 => n_1703, B1 => new_corner_count(28), B2 => n_1704, Z => n_246);
  g30189 : AO22D0BWP7T port map(A1 => n_1677, A2 => n_1703, B1 => new_corner_count(25), B2 => n_1704, Z => n_245);
  g30190 : AO22D0BWP7T port map(A1 => n_1682, A2 => n_1703, B1 => new_corner_count(20), B2 => FE_OFN3_n_1704, Z => n_244);
  g30191 : AO22D0BWP7T port map(A1 => n_1678, A2 => n_1703, B1 => new_corner_count(24), B2 => n_1704, Z => n_243);
  g30192 : AO22D0BWP7T port map(A1 => n_1687, A2 => n_1703, B1 => new_corner_count(15), B2 => FE_OFN3_n_1704, Z => n_242);
  g30193 : AO22D0BWP7T port map(A1 => n_1686, A2 => n_1703, B1 => new_corner_count(16), B2 => FE_OFN3_n_1704, Z => n_241);
  g30194 : NR4D0BWP7T port map(A1 => n_1568, A2 => n_1569, A3 => n_1565, A4 => n_1566, ZN => n_240);
  g30195 : AOI22D0BWP7T port map(A1 => n_152, A2 => snake_output2(5), B1 => N(0), B2 => snake_output3(5), ZN => n_239);
  g30196 : AOI22D0BWP7T port map(A1 => n_153, A2 => snake_output5(5), B1 => N(1), B2 => snake_output7(5), ZN => n_238);
  g30197 : AOI211D0BWP7T port map(A1 => n_1570, A2 => n_1578, B => n_1564, C => n_1567, ZN => n_237);
  g30335 : INVD0BWP7T port map(I => n_228, ZN => n_229);
  g30336 : CKND1BWP7T port map(I => n_225, ZN => n_224);
  g30337 : CKND1BWP7T port map(I => n_217, ZN => n_218);
  g30338 : INVD0BWP7T port map(I => n_214, ZN => n_213);
  g30339 : INVD0BWP7T port map(I => n_212, ZN => n_211);
  g30340 : INVD1BWP7T port map(I => n_208, ZN => n_209);
  g30341 : INVD1BWP7T port map(I => n_206, ZN => n_207);
  g30342 : INVD0BWP7T port map(I => n_205, ZN => n_204);
  g30343 : INVD0BWP7T port map(I => n_203, ZN => n_202);
  g30344 : INVD1BWP7T port map(I => n_195, ZN => n_194);
  g30345 : INVD0BWP7T port map(I => n_193, ZN => n_192);
  g30415 : INR2D0BWP7T port map(A1 => new_N(3), B1 => n_1739, ZN => n_191);
  g30416 : OR2D0BWP7T port map(A1 => n_1739, A2 => new_N(0), Z => n_190);
  g30417 : INR2D0BWP7T port map(A1 => new_N(31), B1 => n_1739, ZN => n_189);
  g30418 : INR2D0BWP7T port map(A1 => new_N(30), B1 => n_1739, ZN => n_188);
  g30419 : NR2D0BWP7T port map(A1 => n_1584, A2 => n_1583, ZN => n_187);
  g30420 : INR2D0BWP7T port map(A1 => new_N(28), B1 => n_1739, ZN => n_186);
  g30421 : INR2D0BWP7T port map(A1 => new_N(27), B1 => n_1739, ZN => n_185);
  g30422 : INR2D0BWP7T port map(A1 => new_N(26), B1 => n_1739, ZN => n_184);
  g30423 : INR2D0BWP7T port map(A1 => new_N(24), B1 => n_1739, ZN => n_183);
  g30424 : INR2D0BWP7T port map(A1 => new_N(29), B1 => n_1739, ZN => n_182);
  g30425 : INR2D0BWP7T port map(A1 => new_N(20), B1 => n_1739, ZN => n_181);
  g30426 : INR2D0BWP7T port map(A1 => new_N(16), B1 => n_1739, ZN => n_180);
  g30427 : INR2D0BWP7T port map(A1 => new_N(19), B1 => n_1739, ZN => n_179);
  g30428 : INR2D0BWP7T port map(A1 => new_N(13), B1 => n_1739, ZN => n_178);
  g30429 : INR2D0BWP7T port map(A1 => new_N(15), B1 => n_1739, ZN => n_177);
  g30430 : INR2D0BWP7T port map(A1 => new_N(18), B1 => n_1739, ZN => n_176);
  g30431 : INR2D0BWP7T port map(A1 => new_N(14), B1 => n_1739, ZN => n_175);
  g30432 : INR2D0BWP7T port map(A1 => new_N(10), B1 => n_1739, ZN => n_174);
  g30433 : INR2D0BWP7T port map(A1 => new_N(7), B1 => n_1739, ZN => n_173);
  g30434 : INR2D0BWP7T port map(A1 => new_N(12), B1 => n_1739, ZN => n_172);
  g30435 : INR2D0BWP7T port map(A1 => new_N(21), B1 => n_1739, ZN => n_171);
  g30436 : INR2D0BWP7T port map(A1 => new_N(6), B1 => n_1739, ZN => n_170);
  g30437 : INR2D0BWP7T port map(A1 => new_N(5), B1 => n_1739, ZN => n_169);
  g30438 : INR2D0BWP7T port map(A1 => new_N(25), B1 => n_1739, ZN => n_168);
  g30439 : INR2D0BWP7T port map(A1 => new_N(11), B1 => n_1739, ZN => n_167);
  g30440 : INR2D0BWP7T port map(A1 => new_N(17), B1 => n_1739, ZN => n_166);
  g30441 : INR2D0BWP7T port map(A1 => new_N(4), B1 => n_1739, ZN => n_165);
  g30442 : ND2D0BWP7T port map(A1 => n_1734, A2 => send_corner_flag, ZN => n_164);
  g30443 : INR2D0BWP7T port map(A1 => new_N(2), B1 => n_1739, ZN => n_163);
  g30444 : INR2D0BWP7T port map(A1 => new_N(1), B1 => n_1739, ZN => n_162);
  g30445 : INR2D0BWP7T port map(A1 => new_N(22), B1 => n_1739, ZN => n_161);
  g30446 : INR2D0BWP7T port map(A1 => new_N(8), B1 => n_1739, ZN => n_160);
  g30447 : INR2D0BWP7T port map(A1 => new_N(9), B1 => n_1739, ZN => n_159);
  g30448 : INR2D0BWP7T port map(A1 => new_N(23), B1 => n_1739, ZN => n_158);
  g30449 : INR2D0BWP7T port map(A1 => n_1654, B1 => n_1650, ZN => n_236);
  g30450 : NR2D0BWP7T port map(A1 => n_1699, A2 => n_1701, ZN => n_235);
  g30451 : NR2D0BWP7T port map(A1 => n_148, A2 => N(3), ZN => n_234);
  g30452 : ND2D0BWP7T port map(A1 => n_1740, A2 => corner_count(1), ZN => n_233);
  g30453 : NR2D0BWP7T port map(A1 => n_1733, A2 => n_1738, ZN => n_232);
  g30454 : NR2D0BWP7T port map(A1 => n_1740, A2 => corner_count(0), ZN => n_231);
  g30455 : ND2D0BWP7T port map(A1 => n_1734, A2 => n_147, ZN => n_230);
  g30456 : NR2D0BWP7T port map(A1 => corner_count(1), A2 => corner_count(2), ZN => n_228);
  g30457 : NR2D0BWP7T port map(A1 => n_1740, A2 => n_146, ZN => n_227);
  g30458 : NR2D0BWP7T port map(A1 => n_148, A2 => N(1), ZN => n_226);
  g30459 : NR2D0BWP7T port map(A1 => n_153, A2 => N(2), ZN => n_225);
  g30460 : NR2D0BWP7T port map(A1 => n_154, A2 => n_149, ZN => n_223);
  g30461 : NR2D0BWP7T port map(A1 => n_1700, A2 => corner_count(0), ZN => n_222);
  g30462 : ND2D0BWP7T port map(A1 => N(2), A2 => N(1), ZN => n_221);
  g30463 : ND2D0BWP7T port map(A1 => n_1700, A2 => n_146, ZN => n_220);
  g30464 : NR2D0BWP7T port map(A1 => N(2), A2 => N(1), ZN => n_219);
  g30465 : ND2D0BWP7T port map(A1 => n_1700, A2 => corner_count(0), ZN => n_217);
  g30466 : ND2D0BWP7T port map(A1 => n_152, A2 => n_153, ZN => n_216);
  g30467 : ND2D0BWP7T port map(A1 => n_148, A2 => n_149, ZN => n_215);
  g30468 : NR2D0BWP7T port map(A1 => n_154, A2 => n_147, ZN => n_214);
  g30469 : NR2D0BWP7T port map(A1 => n_1700, A2 => n_146, ZN => n_212);
  g30470 : ND2D0BWP7T port map(A1 => N(0), A2 => N(1), ZN => n_210);
  g30471 : IND2D0BWP7T port map(A1 => corner_check(5), B1 => n_1653, ZN => n_208);
  g30472 : ND2D0BWP7T port map(A1 => n_1653, A2 => corner_check(5), ZN => n_206);
  g30473 : IND2D0BWP7T port map(A1 => corner_check(5), B1 => n_1732, ZN => n_205);
  g30474 : ND2D0BWP7T port map(A1 => n_1732, A2 => corner_check(5), ZN => n_203);
  g30475 : CKND2D1BWP7T port map(A1 => n_1670, A2 => new_tail(1), ZN => n_201);
  g30476 : CKND2D1BWP7T port map(A1 => n_1670, A2 => new_tail(2), ZN => n_200);
  g30477 : CKND2D1BWP7T port map(A1 => n_1670, A2 => new_tail(0), ZN => n_199);
  g30478 : CKND2D1BWP7T port map(A1 => n_1670, A2 => new_tail(3), ZN => n_198);
  g30479 : CKND2D1BWP7T port map(A1 => n_1670, A2 => new_tail(5), ZN => n_197);
  g30480 : CKND2D1BWP7T port map(A1 => n_1670, A2 => new_tail(4), ZN => n_196);
  g30481 : NR2D0BWP7T port map(A1 => FE_OFN3_n_1704, A2 => n_1739, ZN => n_195);
  g30482 : NR2D1P5BWP7T port map(A1 => n_1732, A2 => n_1653, ZN => n_193);
  g30484 : INVD1BWP7T port map(I => reset, ZN => n_157);
  g30485 : INVD0BWP7T port map(I => n_1701, ZN => n_156);
  g30487 : INVD0BWP7T port map(I => n_1734, ZN => n_154);
  g30488 : INVD0BWP7T port map(I => N(1), ZN => n_153);
  g30489 : INVD0BWP7T port map(I => N(0), ZN => n_152);
  g30490 : INVD1BWP7T port map(I => n_1703, ZN => n_151);
  g30492 : CKND1BWP7T port map(I => n_1700, ZN => n_150);
  g30493 : INVD1BWP7T port map(I => N(3), ZN => n_149);
  g30494 : INVD1BWP7T port map(I => N(2), ZN => n_148);
  g30495 : INVD1BWP7T port map(I => N(4), ZN => n_147);
  g30496 : INVD1BWP7T port map(I => corner_count(0), ZN => n_146);
  drc_bufs30993 : INVD5BWP7T port map(I => n_144, ZN => snake_output4(5));
  drc_bufs30994 : INVD1BWP7T port map(I => n_1167, ZN => n_144);
  drc_bufs31041 : INVD5BWP7T port map(I => n_145, ZN => snake_output23(5));
  drc_bufs31042 : INVD1BWP7T port map(I => n_1053, ZN => n_145);
  g12863 : IND3D1BWP7T port map(A1 => n_610, B1 => n_212, B2 => n_1699, ZN => n_1);
  g31088 : INR3D0BWP7T port map(A1 => n_463, B1 => n_535, B2 => n_429, ZN => n_0);
  g31090 : AO21D0BWP7T port map(A1 => n_1210, A2 => new_corner_flag, B => n_1574, Z => n_1747);
  g31091 : ND3D0BWP7T port map(A1 => n_446, A2 => n_164, A3 => n_240, ZN => n_1748);
  state_reg_0 : DFKCND1BWP7T port map(CN => new_state(0), CP => CTS_6, D => n_157, Q => state(0), QN => n_1205);
  state_reg_2 : DFKCND1BWP7T port map(CN => new_state(2), CP => CTS_6, D => n_157, Q => state(2), QN => n_1204);
  g31096 : IND4D0BWP7T port map(A1 => n_1703, B1 => n_1276, B2 => n_1405, B3 => n_1342, ZN => n_1749);
  inc_add_286_38_g321 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_58, A2 => corner_count(31), B1 => inc_add_286_38_n_58, B2 => corner_count(31), ZN => n_1618);
  inc_add_286_38_g322 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_56, A2 => corner_count(30), B1 => inc_add_286_38_n_56, B2 => corner_count(30), ZN => n_1619);
  inc_add_286_38_g323 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_56, B1 => corner_count(30), ZN => inc_add_286_38_n_58);
  inc_add_286_38_g324 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_54, A2 => corner_count(29), B1 => inc_add_286_38_n_54, B2 => corner_count(29), ZN => n_1620);
  inc_add_286_38_g325 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_54, B1 => corner_count(29), ZN => inc_add_286_38_n_56);
  inc_add_286_38_g326 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_52, A2 => corner_count(28), B1 => inc_add_286_38_n_52, B2 => corner_count(28), ZN => n_1621);
  inc_add_286_38_g327 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_52, B1 => corner_count(28), ZN => inc_add_286_38_n_54);
  inc_add_286_38_g328 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_50, A2 => corner_count(27), B1 => inc_add_286_38_n_50, B2 => corner_count(27), ZN => n_1622);
  inc_add_286_38_g329 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_50, B1 => corner_count(27), ZN => inc_add_286_38_n_52);
  inc_add_286_38_g330 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_48, A2 => corner_count(26), B1 => inc_add_286_38_n_48, B2 => corner_count(26), ZN => n_1623);
  inc_add_286_38_g331 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_48, B1 => corner_count(26), ZN => inc_add_286_38_n_50);
  inc_add_286_38_g332 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_46, A2 => corner_count(25), B1 => inc_add_286_38_n_46, B2 => corner_count(25), ZN => n_1624);
  inc_add_286_38_g333 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_46, B1 => corner_count(25), ZN => inc_add_286_38_n_48);
  inc_add_286_38_g334 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_44, A2 => corner_count(24), B1 => inc_add_286_38_n_44, B2 => corner_count(24), ZN => n_1625);
  inc_add_286_38_g335 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_44, B1 => corner_count(24), ZN => inc_add_286_38_n_46);
  inc_add_286_38_g336 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_42, A2 => corner_count(23), B1 => inc_add_286_38_n_42, B2 => corner_count(23), ZN => n_1626);
  inc_add_286_38_g337 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_42, B1 => corner_count(23), ZN => inc_add_286_38_n_44);
  inc_add_286_38_g338 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_40, A2 => corner_count(22), B1 => inc_add_286_38_n_40, B2 => corner_count(22), ZN => n_1627);
  inc_add_286_38_g339 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_40, B1 => corner_count(22), ZN => inc_add_286_38_n_42);
  inc_add_286_38_g340 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_38, A2 => corner_count(21), B1 => inc_add_286_38_n_38, B2 => corner_count(21), ZN => n_1628);
  inc_add_286_38_g341 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_38, B1 => corner_count(21), ZN => inc_add_286_38_n_40);
  inc_add_286_38_g342 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_36, A2 => corner_count(20), B1 => inc_add_286_38_n_36, B2 => corner_count(20), ZN => n_1629);
  inc_add_286_38_g343 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_36, B1 => corner_count(20), ZN => inc_add_286_38_n_38);
  inc_add_286_38_g344 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_34, A2 => corner_count(19), B1 => inc_add_286_38_n_34, B2 => corner_count(19), ZN => n_1630);
  inc_add_286_38_g345 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_34, B1 => corner_count(19), ZN => inc_add_286_38_n_36);
  inc_add_286_38_g346 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_32, A2 => corner_count(18), B1 => inc_add_286_38_n_32, B2 => corner_count(18), ZN => n_1631);
  inc_add_286_38_g347 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_32, B1 => corner_count(18), ZN => inc_add_286_38_n_34);
  inc_add_286_38_g348 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_30, A2 => corner_count(17), B1 => inc_add_286_38_n_30, B2 => corner_count(17), ZN => n_1632);
  inc_add_286_38_g349 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_30, B1 => corner_count(17), ZN => inc_add_286_38_n_32);
  inc_add_286_38_g350 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_28, A2 => corner_count(16), B1 => inc_add_286_38_n_28, B2 => corner_count(16), ZN => n_1633);
  inc_add_286_38_g351 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_28, B1 => corner_count(16), ZN => inc_add_286_38_n_30);
  inc_add_286_38_g352 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_26, A2 => corner_count(15), B1 => inc_add_286_38_n_26, B2 => corner_count(15), ZN => n_1634);
  inc_add_286_38_g353 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_26, B1 => corner_count(15), ZN => inc_add_286_38_n_28);
  inc_add_286_38_g354 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_24, A2 => corner_count(14), B1 => inc_add_286_38_n_24, B2 => corner_count(14), ZN => n_1635);
  inc_add_286_38_g355 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_24, B1 => corner_count(14), ZN => inc_add_286_38_n_26);
  inc_add_286_38_g356 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_22, A2 => corner_count(13), B1 => inc_add_286_38_n_22, B2 => corner_count(13), ZN => n_1636);
  inc_add_286_38_g357 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_22, B1 => corner_count(13), ZN => inc_add_286_38_n_24);
  inc_add_286_38_g358 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_20, A2 => corner_count(12), B1 => inc_add_286_38_n_20, B2 => corner_count(12), ZN => n_1637);
  inc_add_286_38_g359 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_20, B1 => corner_count(12), ZN => inc_add_286_38_n_22);
  inc_add_286_38_g360 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_18, A2 => corner_count(11), B1 => inc_add_286_38_n_18, B2 => corner_count(11), ZN => n_1638);
  inc_add_286_38_g361 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_18, B1 => corner_count(11), ZN => inc_add_286_38_n_20);
  inc_add_286_38_g362 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_16, A2 => corner_count(10), B1 => inc_add_286_38_n_16, B2 => corner_count(10), ZN => n_1639);
  inc_add_286_38_g363 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_16, B1 => corner_count(10), ZN => inc_add_286_38_n_18);
  inc_add_286_38_g364 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_14, A2 => corner_count(9), B1 => inc_add_286_38_n_14, B2 => corner_count(9), ZN => n_1640);
  inc_add_286_38_g365 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_14, B1 => corner_count(9), ZN => inc_add_286_38_n_16);
  inc_add_286_38_g366 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_12, A2 => corner_count(8), B1 => inc_add_286_38_n_12, B2 => corner_count(8), ZN => n_1641);
  inc_add_286_38_g367 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_12, B1 => corner_count(8), ZN => inc_add_286_38_n_14);
  inc_add_286_38_g368 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_10, A2 => corner_count(7), B1 => inc_add_286_38_n_10, B2 => corner_count(7), ZN => n_1642);
  inc_add_286_38_g369 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_10, B1 => corner_count(7), ZN => inc_add_286_38_n_12);
  inc_add_286_38_g370 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_8, A2 => corner_count(6), B1 => inc_add_286_38_n_8, B2 => corner_count(6), ZN => n_1643);
  inc_add_286_38_g371 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_8, B1 => corner_count(6), ZN => inc_add_286_38_n_10);
  inc_add_286_38_g372 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_6, A2 => corner_count(5), B1 => inc_add_286_38_n_6, B2 => corner_count(5), ZN => n_1644);
  inc_add_286_38_g373 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_6, B1 => corner_count(5), ZN => inc_add_286_38_n_8);
  inc_add_286_38_g374 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_4, A2 => corner_count(4), B1 => inc_add_286_38_n_4, B2 => corner_count(4), ZN => n_1645);
  inc_add_286_38_g375 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_4, B1 => corner_count(4), ZN => inc_add_286_38_n_6);
  inc_add_286_38_g376 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_2, A2 => corner_count(3), B1 => inc_add_286_38_n_2, B2 => corner_count(3), ZN => n_1646);
  inc_add_286_38_g377 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_2, B1 => corner_count(3), ZN => inc_add_286_38_n_4);
  inc_add_286_38_g378 : MOAI22D0BWP7T port map(A1 => inc_add_286_38_n_0, A2 => corner_count(2), B1 => inc_add_286_38_n_0, B2 => corner_count(2), ZN => n_1647);
  inc_add_286_38_g379 : IND2D0BWP7T port map(A1 => inc_add_286_38_n_0, B1 => corner_count(2), ZN => inc_add_286_38_n_2);
  inc_add_286_38_g380 : CKXOR2D0BWP7T port map(A1 => corner_count(0), A2 => corner_count(1), Z => n_1648);
  inc_add_286_38_g381 : ND2D0BWP7T port map(A1 => corner_count(0), A2 => corner_count(1), ZN => inc_add_286_38_n_0);
  inc_add_1070_17_g321 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_58, A2 => N(31), B1 => inc_add_1070_17_n_58, B2 => N(31), ZN => n_1587);
  inc_add_1070_17_g322 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_56, A2 => N(30), B1 => inc_add_1070_17_n_56, B2 => N(30), ZN => n_1588);
  inc_add_1070_17_g323 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_56, B1 => N(30), ZN => inc_add_1070_17_n_58);
  inc_add_1070_17_g324 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_54, A2 => N(29), B1 => inc_add_1070_17_n_54, B2 => N(29), ZN => n_1589);
  inc_add_1070_17_g325 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_54, B1 => N(29), ZN => inc_add_1070_17_n_56);
  inc_add_1070_17_g326 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_52, A2 => N(28), B1 => inc_add_1070_17_n_52, B2 => N(28), ZN => n_1590);
  inc_add_1070_17_g327 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_52, B1 => N(28), ZN => inc_add_1070_17_n_54);
  inc_add_1070_17_g328 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_50, A2 => N(27), B1 => inc_add_1070_17_n_50, B2 => N(27), ZN => n_1591);
  inc_add_1070_17_g329 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_50, B1 => N(27), ZN => inc_add_1070_17_n_52);
  inc_add_1070_17_g330 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_48, A2 => N(26), B1 => inc_add_1070_17_n_48, B2 => N(26), ZN => n_1592);
  inc_add_1070_17_g331 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_48, B1 => N(26), ZN => inc_add_1070_17_n_50);
  inc_add_1070_17_g332 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_46, A2 => N(25), B1 => inc_add_1070_17_n_46, B2 => N(25), ZN => n_1593);
  inc_add_1070_17_g333 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_46, B1 => N(25), ZN => inc_add_1070_17_n_48);
  inc_add_1070_17_g334 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_44, A2 => N(24), B1 => inc_add_1070_17_n_44, B2 => N(24), ZN => n_1594);
  inc_add_1070_17_g335 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_44, B1 => N(24), ZN => inc_add_1070_17_n_46);
  inc_add_1070_17_g336 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_42, A2 => N(23), B1 => inc_add_1070_17_n_42, B2 => N(23), ZN => n_1595);
  inc_add_1070_17_g337 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_42, B1 => N(23), ZN => inc_add_1070_17_n_44);
  inc_add_1070_17_g338 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_40, A2 => N(22), B1 => inc_add_1070_17_n_40, B2 => N(22), ZN => n_1596);
  inc_add_1070_17_g339 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_40, B1 => N(22), ZN => inc_add_1070_17_n_42);
  inc_add_1070_17_g340 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_38, A2 => N(21), B1 => inc_add_1070_17_n_38, B2 => N(21), ZN => n_1597);
  inc_add_1070_17_g341 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_38, B1 => N(21), ZN => inc_add_1070_17_n_40);
  inc_add_1070_17_g342 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_36, A2 => N(20), B1 => inc_add_1070_17_n_36, B2 => N(20), ZN => n_1598);
  inc_add_1070_17_g343 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_36, B1 => N(20), ZN => inc_add_1070_17_n_38);
  inc_add_1070_17_g344 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_34, A2 => N(19), B1 => inc_add_1070_17_n_34, B2 => N(19), ZN => n_1599);
  inc_add_1070_17_g345 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_34, B1 => N(19), ZN => inc_add_1070_17_n_36);
  inc_add_1070_17_g346 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_32, A2 => N(18), B1 => inc_add_1070_17_n_32, B2 => N(18), ZN => n_1600);
  inc_add_1070_17_g347 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_32, B1 => N(18), ZN => inc_add_1070_17_n_34);
  inc_add_1070_17_g348 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_30, A2 => N(17), B1 => inc_add_1070_17_n_30, B2 => N(17), ZN => n_1601);
  inc_add_1070_17_g349 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_30, B1 => N(17), ZN => inc_add_1070_17_n_32);
  inc_add_1070_17_g350 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_28, A2 => N(16), B1 => inc_add_1070_17_n_28, B2 => N(16), ZN => n_1602);
  inc_add_1070_17_g351 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_28, B1 => N(16), ZN => inc_add_1070_17_n_30);
  inc_add_1070_17_g352 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_26, A2 => N(15), B1 => inc_add_1070_17_n_26, B2 => N(15), ZN => n_1603);
  inc_add_1070_17_g353 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_26, B1 => N(15), ZN => inc_add_1070_17_n_28);
  inc_add_1070_17_g354 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_24, A2 => N(14), B1 => inc_add_1070_17_n_24, B2 => N(14), ZN => n_1604);
  inc_add_1070_17_g355 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_24, B1 => N(14), ZN => inc_add_1070_17_n_26);
  inc_add_1070_17_g356 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_22, A2 => N(13), B1 => inc_add_1070_17_n_22, B2 => N(13), ZN => n_1605);
  inc_add_1070_17_g357 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_22, B1 => N(13), ZN => inc_add_1070_17_n_24);
  inc_add_1070_17_g358 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_20, A2 => N(12), B1 => inc_add_1070_17_n_20, B2 => N(12), ZN => n_1606);
  inc_add_1070_17_g359 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_20, B1 => N(12), ZN => inc_add_1070_17_n_22);
  inc_add_1070_17_g360 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_18, A2 => N(11), B1 => inc_add_1070_17_n_18, B2 => N(11), ZN => n_1607);
  inc_add_1070_17_g361 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_18, B1 => N(11), ZN => inc_add_1070_17_n_20);
  inc_add_1070_17_g362 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_16, A2 => N(10), B1 => inc_add_1070_17_n_16, B2 => N(10), ZN => n_1608);
  inc_add_1070_17_g363 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_16, B1 => N(10), ZN => inc_add_1070_17_n_18);
  inc_add_1070_17_g364 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_14, A2 => N(9), B1 => inc_add_1070_17_n_14, B2 => N(9), ZN => n_1609);
  inc_add_1070_17_g365 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_14, B1 => N(9), ZN => inc_add_1070_17_n_16);
  inc_add_1070_17_g366 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_12, A2 => N(8), B1 => inc_add_1070_17_n_12, B2 => N(8), ZN => n_1610);
  inc_add_1070_17_g367 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_12, B1 => N(8), ZN => inc_add_1070_17_n_14);
  inc_add_1070_17_g368 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_10, A2 => N(7), B1 => inc_add_1070_17_n_10, B2 => N(7), ZN => n_1611);
  inc_add_1070_17_g369 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_10, B1 => N(7), ZN => inc_add_1070_17_n_12);
  inc_add_1070_17_g370 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_8, A2 => N(6), B1 => inc_add_1070_17_n_8, B2 => N(6), ZN => n_1612);
  inc_add_1070_17_g371 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_8, B1 => N(6), ZN => inc_add_1070_17_n_10);
  inc_add_1070_17_g372 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_6, A2 => N(5), B1 => inc_add_1070_17_n_6, B2 => N(5), ZN => n_1613);
  inc_add_1070_17_g373 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_6, B1 => N(5), ZN => inc_add_1070_17_n_8);
  inc_add_1070_17_g374 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_4, A2 => N(4), B1 => inc_add_1070_17_n_4, B2 => N(4), ZN => n_1614);
  inc_add_1070_17_g375 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_4, B1 => N(4), ZN => inc_add_1070_17_n_6);
  inc_add_1070_17_g376 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_2, A2 => N(3), B1 => inc_add_1070_17_n_2, B2 => N(3), ZN => n_1615);
  inc_add_1070_17_g377 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_2, B1 => N(3), ZN => inc_add_1070_17_n_4);
  inc_add_1070_17_g378 : MOAI22D0BWP7T port map(A1 => inc_add_1070_17_n_0, A2 => N(2), B1 => inc_add_1070_17_n_0, B2 => N(2), ZN => n_1616);
  inc_add_1070_17_g379 : IND2D0BWP7T port map(A1 => inc_add_1070_17_n_0, B1 => N(2), ZN => inc_add_1070_17_n_2);
  inc_add_1070_17_g380 : CKXOR2D0BWP7T port map(A1 => N(0), A2 => N(1), Z => n_1617);
  inc_add_1070_17_g381 : ND2D0BWP7T port map(A1 => N(0), A2 => N(1), ZN => inc_add_1070_17_n_0);
  sub_868_22_g709 : MOAI22D0BWP7T port map(A1 => sub_868_22_n_58, A2 => corner_count(31), B1 => sub_868_22_n_58, B2 => corner_count(31), ZN => n_1671);
  sub_868_22_g710 : IOA21D0BWP7T port map(A1 => sub_868_22_n_56, A2 => corner_count(30), B => sub_868_22_n_58, ZN => n_1672);
  sub_868_22_g711 : OR2D0BWP7T port map(A1 => sub_868_22_n_56, A2 => corner_count(30), Z => sub_868_22_n_58);
  sub_868_22_g712 : IOA21D0BWP7T port map(A1 => sub_868_22_n_54, A2 => corner_count(29), B => sub_868_22_n_56, ZN => n_1673);
  sub_868_22_g713 : OR2D0BWP7T port map(A1 => sub_868_22_n_54, A2 => corner_count(29), Z => sub_868_22_n_56);
  sub_868_22_g714 : IOA21D0BWP7T port map(A1 => sub_868_22_n_52, A2 => corner_count(28), B => sub_868_22_n_54, ZN => n_1674);
  sub_868_22_g715 : OR2D0BWP7T port map(A1 => sub_868_22_n_52, A2 => corner_count(28), Z => sub_868_22_n_54);
  sub_868_22_g716 : IOA21D0BWP7T port map(A1 => sub_868_22_n_50, A2 => corner_count(27), B => sub_868_22_n_52, ZN => n_1675);
  sub_868_22_g717 : OR2D0BWP7T port map(A1 => sub_868_22_n_50, A2 => corner_count(27), Z => sub_868_22_n_52);
  sub_868_22_g718 : IOA21D0BWP7T port map(A1 => sub_868_22_n_48, A2 => corner_count(26), B => sub_868_22_n_50, ZN => n_1676);
  sub_868_22_g719 : OR2D0BWP7T port map(A1 => sub_868_22_n_48, A2 => corner_count(26), Z => sub_868_22_n_50);
  sub_868_22_g720 : IOA21D0BWP7T port map(A1 => sub_868_22_n_46, A2 => corner_count(25), B => sub_868_22_n_48, ZN => n_1677);
  sub_868_22_g721 : OR2D0BWP7T port map(A1 => sub_868_22_n_46, A2 => corner_count(25), Z => sub_868_22_n_48);
  sub_868_22_g722 : IOA21D0BWP7T port map(A1 => sub_868_22_n_44, A2 => corner_count(24), B => sub_868_22_n_46, ZN => n_1678);
  sub_868_22_g723 : OR2D0BWP7T port map(A1 => sub_868_22_n_44, A2 => corner_count(24), Z => sub_868_22_n_46);
  sub_868_22_g724 : IOA21D0BWP7T port map(A1 => sub_868_22_n_42, A2 => corner_count(23), B => sub_868_22_n_44, ZN => n_1679);
  sub_868_22_g725 : OR2D0BWP7T port map(A1 => sub_868_22_n_42, A2 => corner_count(23), Z => sub_868_22_n_44);
  sub_868_22_g726 : IOA21D0BWP7T port map(A1 => sub_868_22_n_40, A2 => corner_count(22), B => sub_868_22_n_42, ZN => n_1680);
  sub_868_22_g727 : OR2D0BWP7T port map(A1 => sub_868_22_n_40, A2 => corner_count(22), Z => sub_868_22_n_42);
  sub_868_22_g728 : IOA21D0BWP7T port map(A1 => sub_868_22_n_38, A2 => corner_count(21), B => sub_868_22_n_40, ZN => n_1681);
  sub_868_22_g729 : OR2D0BWP7T port map(A1 => sub_868_22_n_38, A2 => corner_count(21), Z => sub_868_22_n_40);
  sub_868_22_g730 : IOA21D0BWP7T port map(A1 => sub_868_22_n_36, A2 => corner_count(20), B => sub_868_22_n_38, ZN => n_1682);
  sub_868_22_g731 : OR2D0BWP7T port map(A1 => sub_868_22_n_36, A2 => corner_count(20), Z => sub_868_22_n_38);
  sub_868_22_g732 : IOA21D0BWP7T port map(A1 => sub_868_22_n_34, A2 => corner_count(19), B => sub_868_22_n_36, ZN => n_1683);
  sub_868_22_g733 : OR2D0BWP7T port map(A1 => sub_868_22_n_34, A2 => corner_count(19), Z => sub_868_22_n_36);
  sub_868_22_g734 : IOA21D0BWP7T port map(A1 => sub_868_22_n_32, A2 => corner_count(18), B => sub_868_22_n_34, ZN => n_1684);
  sub_868_22_g735 : OR2D0BWP7T port map(A1 => sub_868_22_n_32, A2 => corner_count(18), Z => sub_868_22_n_34);
  sub_868_22_g736 : IOA21D0BWP7T port map(A1 => sub_868_22_n_30, A2 => corner_count(17), B => sub_868_22_n_32, ZN => n_1685);
  sub_868_22_g737 : OR2D0BWP7T port map(A1 => sub_868_22_n_30, A2 => corner_count(17), Z => sub_868_22_n_32);
  sub_868_22_g738 : IOA21D0BWP7T port map(A1 => sub_868_22_n_28, A2 => corner_count(16), B => sub_868_22_n_30, ZN => n_1686);
  sub_868_22_g739 : OR2D0BWP7T port map(A1 => sub_868_22_n_28, A2 => corner_count(16), Z => sub_868_22_n_30);
  sub_868_22_g740 : IOA21D0BWP7T port map(A1 => sub_868_22_n_26, A2 => corner_count(15), B => sub_868_22_n_28, ZN => n_1687);
  sub_868_22_g741 : OR2D0BWP7T port map(A1 => sub_868_22_n_26, A2 => corner_count(15), Z => sub_868_22_n_28);
  sub_868_22_g742 : IOA21D0BWP7T port map(A1 => sub_868_22_n_24, A2 => corner_count(14), B => sub_868_22_n_26, ZN => n_1688);
  sub_868_22_g743 : OR2D0BWP7T port map(A1 => sub_868_22_n_24, A2 => corner_count(14), Z => sub_868_22_n_26);
  sub_868_22_g744 : IOA21D0BWP7T port map(A1 => sub_868_22_n_22, A2 => corner_count(13), B => sub_868_22_n_24, ZN => n_1689);
  sub_868_22_g745 : OR2D0BWP7T port map(A1 => sub_868_22_n_22, A2 => corner_count(13), Z => sub_868_22_n_24);
  sub_868_22_g746 : IOA21D0BWP7T port map(A1 => sub_868_22_n_20, A2 => corner_count(12), B => sub_868_22_n_22, ZN => n_1690);
  sub_868_22_g747 : OR2D0BWP7T port map(A1 => sub_868_22_n_20, A2 => corner_count(12), Z => sub_868_22_n_22);
  sub_868_22_g748 : IOA21D0BWP7T port map(A1 => sub_868_22_n_18, A2 => corner_count(11), B => sub_868_22_n_20, ZN => n_1691);
  sub_868_22_g749 : OR2D0BWP7T port map(A1 => sub_868_22_n_18, A2 => corner_count(11), Z => sub_868_22_n_20);
  sub_868_22_g750 : IOA21D0BWP7T port map(A1 => sub_868_22_n_16, A2 => corner_count(10), B => sub_868_22_n_18, ZN => n_1692);
  sub_868_22_g751 : OR2D0BWP7T port map(A1 => sub_868_22_n_16, A2 => corner_count(10), Z => sub_868_22_n_18);
  sub_868_22_g752 : IOA21D0BWP7T port map(A1 => sub_868_22_n_14, A2 => corner_count(9), B => sub_868_22_n_16, ZN => n_1693);
  sub_868_22_g753 : OR2D0BWP7T port map(A1 => sub_868_22_n_14, A2 => corner_count(9), Z => sub_868_22_n_16);
  sub_868_22_g754 : IOA21D0BWP7T port map(A1 => sub_868_22_n_12, A2 => corner_count(8), B => sub_868_22_n_14, ZN => n_1694);
  sub_868_22_g755 : OR2D0BWP7T port map(A1 => sub_868_22_n_12, A2 => corner_count(8), Z => sub_868_22_n_14);
  sub_868_22_g756 : IOA21D0BWP7T port map(A1 => sub_868_22_n_10, A2 => corner_count(7), B => sub_868_22_n_12, ZN => n_1695);
  sub_868_22_g757 : OR2D0BWP7T port map(A1 => sub_868_22_n_10, A2 => corner_count(7), Z => sub_868_22_n_12);
  sub_868_22_g758 : IOA21D0BWP7T port map(A1 => sub_868_22_n_8, A2 => corner_count(6), B => sub_868_22_n_10, ZN => n_1696);
  sub_868_22_g759 : OR2D0BWP7T port map(A1 => sub_868_22_n_8, A2 => corner_count(6), Z => sub_868_22_n_10);
  sub_868_22_g760 : IOA21D0BWP7T port map(A1 => sub_868_22_n_6, A2 => corner_count(5), B => sub_868_22_n_8, ZN => n_1697);
  sub_868_22_g761 : OR2D0BWP7T port map(A1 => sub_868_22_n_6, A2 => corner_count(5), Z => sub_868_22_n_8);
  sub_868_22_g762 : IOA21D0BWP7T port map(A1 => sub_868_22_n_4, A2 => corner_count(4), B => sub_868_22_n_6, ZN => n_1698);
  sub_868_22_g763 : OR2D0BWP7T port map(A1 => sub_868_22_n_4, A2 => corner_count(4), Z => sub_868_22_n_6);
  sub_868_22_g764 : IOA21D0BWP7T port map(A1 => sub_868_22_n_2, A2 => corner_count(3), B => sub_868_22_n_4, ZN => n_1699);
  sub_868_22_g765 : OR2D0BWP7T port map(A1 => sub_868_22_n_2, A2 => corner_count(3), Z => sub_868_22_n_4);
  sub_868_22_g766 : IOA21D0BWP7T port map(A1 => sub_868_22_n_0, A2 => corner_count(2), B => sub_868_22_n_2, ZN => n_1700);
  sub_868_22_g767 : OR2D0BWP7T port map(A1 => sub_868_22_n_0, A2 => corner_count(2), Z => sub_868_22_n_2);
  sub_868_22_g768 : IOA21D0BWP7T port map(A1 => corner_count(1), A2 => corner_count(0), B => sub_868_22_n_0, ZN => n_1701);
  sub_868_22_g769 : OR2D0BWP7T port map(A1 => corner_count(0), A2 => corner_count(1), Z => sub_868_22_n_0);
  tie_0_cell : TIELBWP7T port map(ZN => FE_OFN5_audio_0);

end routed;
