configuration shift_register_behaviour_cfg of shift_register is
   for behaviour
   end for;
end shift_register_behaviour_cfg;
