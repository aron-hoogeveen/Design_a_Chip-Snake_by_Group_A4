configuration itemgenerator_tb_behaviour_cfg of itemgenerator_tb is
   for behaviour
      for all: itemgenerator use configuration work.itemgenerator_behaviour_cfg;
      end for;
   end for;
end itemgenerator_tb_behaviour_cfg;
