library IEEE;
use IEEE.std_logic_1164.ALL;

entity image_gen_tb is
end image_gen_tb;

